// file: ibert_7series_gtx_0.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series 
//  /   /         Filename : example_ibert_7series_gtx_0
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module example_ibert_7series_gtx_0
// Generated by Xilinx IBERT_7S 
//////////////////////////////////////////////////////////////////////////////


`define C_NUM_QUADS 1
`define C_REFCLKS_USED 1
module example_ibert_7series_gtx_0
(
  // GT top level ports
  output [(4*`C_NUM_QUADS)-1:0]		TXN_O,
  output [(4*`C_NUM_QUADS)-1:0]		TXP_O,
  input  [(4*`C_NUM_QUADS)-1:0]    	RXN_I,
  input  [(4*`C_NUM_QUADS)-1:0]   	RXP_I,
  input  [`C_REFCLKS_USED-1:0]        	GTREFCLK0P_I,
  input  [`C_REFCLKS_USED-1:0]        	GTREFCLK0N_I,
  input  [`C_REFCLKS_USED-1:0]        	GTREFCLK1P_I,
  input  [`C_REFCLKS_USED-1:0]        	GTREFCLK1N_I,
  output SFP1_TX_DIS,
  output SFP2_TX_DIS
);

  //
  // Ibert refclk internal signals
  //
  wire   [`C_NUM_QUADS-1:0]        	gtrefclk0_i;
  wire   [`C_NUM_QUADS-1:0]        	gtrefclk1_i;
  wire   [`C_REFCLKS_USED-1:0]        	refclk0_i;
  wire   [`C_REFCLKS_USED-1:0]        	refclk1_i;

  //
  // Refclk IBUFDS instantiations
  //

    IBUFDS_GTE2 u_buf_q1_clk1
      (
        .O            (refclk1_i[0]),
        .ODIV2        (),
        .CEB          (1'b0),
        .I            (GTREFCLK1P_I[0]),
        .IB           (GTREFCLK1N_I[0])
      );

  //
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gtrefclk0_i[0] = 1'b0;
  assign gtrefclk1_i[0] = refclk1_i[0];





  //
  // IBERT core instantiation
  //
  ibert_7series_gtx_0 u_ibert_core
    (
      .TXN_O(TXN_O),
      .TXP_O(TXP_O),
      .RXN_I(RXN_I),
      .RXP_I(RXP_I),
      .GTREFCLK0_I(gtrefclk0_i),
      .GTREFCLK1_I(gtrefclk1_i)
    );

// The finisar FTLF8524P2BNV fibre channel SFP transceiver datasheet
// https://edt.com/wp-content/uploads/2018/06/FTLF8524P2BNV.pdf
// says the " Laser output disabled on high or open" for the Tdis pin
// The TOSING_160T schematic shows the TX_DIS signals has a 4.7K pull-up to 3.3V.
// Therefore, need to drive these signals low to enable the laser.
assign SFP1_TX_DIS = 0;
assign SFP2_TX_DIS = 0;

endmodule

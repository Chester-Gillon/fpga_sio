-- vim: ts=4 sw=4 expandtab

-- THIS IS GENERATED VHDL CODE.
-- https://bues.ch/h/crcgen
-- 
-- This code is Public Domain.
-- Permission to use, copy, modify, and/or distribute this software for any
-- purpose with or without fee is hereby granted.
-- 
-- THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
-- WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
-- MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR ANY
-- SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES WHATSOEVER
-- RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN ACTION OF CONTRACT,
-- NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF OR IN CONNECTION WITH THE
-- USE OR PERFORMANCE OF THIS SOFTWARE.

-- CRC polynomial coefficients: x^64 + x^62 + x^57 + x^55 + x^54 + x^53 + x^52 + x^47 + x^46 + x^45 + x^40 + x^39 + x^38 + x^37 + x^35 + x^33 + x^32 + x^31 + x^29 + x^27 + x^24 + x^23 + x^22 + x^21 + x^19 + x^17 + x^13 + x^12 + x^10 + x^9 + x^7 + x^4 + x + 1
--                              0xC96C5795D7870F42 (hex)
-- CRC width:                   64 bits
-- CRC shift direction:         right (little endian)
-- Input word width:            512 bits

library IEEE;
use IEEE.std_logic_1164.all;

entity crc is
    port (
        crc_in: in std_logic_vector(63 downto 0);
        data_in: in std_logic_vector(511 downto 0);
        crc_out: out std_logic_vector(63 downto 0)
    );
end entity crc;

architecture Behavioral of crc is
begin
    crc_out(0) <= crc_in(0) xor crc_in(2) xor crc_in(5) xor crc_in(7) xor crc_in(8) xor crc_in(10) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(21) xor crc_in(22) xor crc_in(24) xor crc_in(32) xor crc_in(36) xor crc_in(41) xor crc_in(43) xor crc_in(45) xor crc_in(47) xor crc_in(50) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(58) xor crc_in(59) xor crc_in(62) xor data_in(0) xor data_in(2) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(21) xor data_in(22) xor data_in(24) xor data_in(32) xor data_in(36) xor data_in(41) xor data_in(43) xor data_in(45) xor data_in(47) xor data_in(50) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(58) xor data_in(59) xor data_in(62) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(74) xor data_in(76) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(82) xor data_in(83) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(92) xor data_in(95) xor data_in(102) xor data_in(103) xor data_in(104) xor data_in(108) xor data_in(110) xor data_in(111) xor data_in(113) xor data_in(114) xor data_in(119) xor data_in(120) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(126) xor data_in(129) xor data_in(130) xor data_in(132) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(142) xor data_in(143) xor data_in(146) xor data_in(150) xor data_in(151) xor data_in(152) xor data_in(154) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(158) xor data_in(160) xor data_in(164) xor data_in(165) xor data_in(166) xor data_in(167) xor data_in(168) xor data_in(170) xor data_in(171) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(181) xor data_in(182) xor data_in(184) xor data_in(186) xor data_in(190) xor data_in(194) xor data_in(197) xor data_in(200) xor data_in(204) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(208) xor data_in(211) xor data_in(212) xor data_in(214) xor data_in(216) xor data_in(218) xor data_in(223) xor data_in(224) xor data_in(225) xor data_in(226) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(239) xor data_in(242) xor data_in(245) xor data_in(252) xor data_in(254) xor data_in(258) xor data_in(262) xor data_in(263) xor data_in(264) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(275) xor data_in(276) xor data_in(278) xor data_in(281) xor data_in(287) xor data_in(288) xor data_in(291) xor data_in(295) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(302) xor data_in(303) xor data_in(304) xor data_in(309) xor data_in(313) xor data_in(314) xor data_in(318) xor data_in(320) xor data_in(323) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(338) xor data_in(339) xor data_in(340) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(348) xor data_in(349) xor data_in(352) xor data_in(353) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(362) xor data_in(363) xor data_in(364) xor data_in(367) xor data_in(368) xor data_in(372) xor data_in(373) xor data_in(379) xor data_in(380) xor data_in(382) xor data_in(385) xor data_in(387) xor data_in(388) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(395) xor data_in(397) xor data_in(398) xor data_in(400) xor data_in(405) xor data_in(408) xor data_in(409) xor data_in(412) xor data_in(413) xor data_in(416) xor data_in(417) xor data_in(419) xor data_in(420) xor data_in(421) xor data_in(423) xor data_in(424) xor data_in(429) xor data_in(430) xor data_in(431) xor data_in(434) xor data_in(435) xor data_in(438) xor data_in(439) xor data_in(442) xor data_in(449) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(463) xor data_in(466) xor data_in(470) xor data_in(471) xor data_in(474) xor data_in(475) xor data_in(477) xor data_in(478) xor data_in(484) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(491) xor data_in(493) xor data_in(496) xor data_in(498) xor data_in(499) xor data_in(503) xor data_in(504) xor data_in(505) xor data_in(506) xor data_in(508) xor data_in(510);
    crc_out(1) <= crc_in(0) xor crc_in(1) xor crc_in(3) xor crc_in(6) xor crc_in(8) xor crc_in(9) xor crc_in(11) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(22) xor crc_in(23) xor crc_in(25) xor crc_in(33) xor crc_in(37) xor crc_in(42) xor crc_in(44) xor crc_in(46) xor crc_in(48) xor crc_in(51) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(59) xor crc_in(60) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(6) xor data_in(8) xor data_in(9) xor data_in(11) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(22) xor data_in(23) xor data_in(25) xor data_in(33) xor data_in(37) xor data_in(42) xor data_in(44) xor data_in(46) xor data_in(48) xor data_in(51) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(59) xor data_in(60) xor data_in(63) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(75) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(83) xor data_in(84) xor data_in(86) xor data_in(87) xor data_in(88) xor data_in(93) xor data_in(96) xor data_in(103) xor data_in(104) xor data_in(105) xor data_in(109) xor data_in(111) xor data_in(112) xor data_in(114) xor data_in(115) xor data_in(120) xor data_in(121) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(127) xor data_in(130) xor data_in(131) xor data_in(133) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(142) xor data_in(143) xor data_in(144) xor data_in(147) xor data_in(151) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(158) xor data_in(159) xor data_in(161) xor data_in(165) xor data_in(166) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(171) xor data_in(172) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(182) xor data_in(183) xor data_in(185) xor data_in(187) xor data_in(191) xor data_in(195) xor data_in(198) xor data_in(201) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(208) xor data_in(209) xor data_in(212) xor data_in(213) xor data_in(215) xor data_in(217) xor data_in(219) xor data_in(224) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(240) xor data_in(243) xor data_in(246) xor data_in(253) xor data_in(255) xor data_in(259) xor data_in(263) xor data_in(264) xor data_in(265) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(270) xor data_in(276) xor data_in(277) xor data_in(279) xor data_in(282) xor data_in(288) xor data_in(289) xor data_in(292) xor data_in(296) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(303) xor data_in(304) xor data_in(305) xor data_in(310) xor data_in(314) xor data_in(315) xor data_in(319) xor data_in(321) xor data_in(324) xor data_in(326) xor data_in(327) xor data_in(328) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(339) xor data_in(340) xor data_in(341) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(349) xor data_in(350) xor data_in(353) xor data_in(354) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(368) xor data_in(369) xor data_in(373) xor data_in(374) xor data_in(380) xor data_in(381) xor data_in(383) xor data_in(386) xor data_in(388) xor data_in(389) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(396) xor data_in(398) xor data_in(399) xor data_in(401) xor data_in(406) xor data_in(409) xor data_in(410) xor data_in(413) xor data_in(414) xor data_in(417) xor data_in(418) xor data_in(420) xor data_in(421) xor data_in(422) xor data_in(424) xor data_in(425) xor data_in(430) xor data_in(431) xor data_in(432) xor data_in(435) xor data_in(436) xor data_in(439) xor data_in(440) xor data_in(443) xor data_in(450) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(463) xor data_in(464) xor data_in(467) xor data_in(471) xor data_in(472) xor data_in(475) xor data_in(476) xor data_in(478) xor data_in(479) xor data_in(485) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(492) xor data_in(494) xor data_in(497) xor data_in(499) xor data_in(500) xor data_in(504) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(509) xor data_in(511);
    crc_out(2) <= crc_in(1) xor crc_in(4) xor crc_in(5) xor crc_in(8) xor crc_in(9) xor crc_in(13) xor crc_in(16) xor crc_in(17) xor crc_in(21) xor crc_in(22) xor crc_in(23) xor crc_in(26) xor crc_in(32) xor crc_in(34) xor crc_in(36) xor crc_in(38) xor crc_in(41) xor crc_in(49) xor crc_in(50) xor crc_in(53) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor data_in(1) xor data_in(4) xor data_in(5) xor data_in(8) xor data_in(9) xor data_in(13) xor data_in(16) xor data_in(17) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(26) xor data_in(32) xor data_in(34) xor data_in(36) xor data_in(38) xor data_in(41) xor data_in(49) xor data_in(50) xor data_in(53) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(64) xor data_in(69) xor data_in(70) xor data_in(73) xor data_in(77) xor data_in(81) xor data_in(83) xor data_in(84) xor data_in(86) xor data_in(88) xor data_in(89) xor data_in(92) xor data_in(94) xor data_in(95) xor data_in(97) xor data_in(102) xor data_in(103) xor data_in(105) xor data_in(106) xor data_in(108) xor data_in(111) xor data_in(112) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(123) xor data_in(125) xor data_in(128) xor data_in(129) xor data_in(130) xor data_in(131) xor data_in(134) xor data_in(136) xor data_in(137) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(148) xor data_in(150) xor data_in(151) xor data_in(153) xor data_in(155) xor data_in(159) xor data_in(162) xor data_in(164) xor data_in(165) xor data_in(169) xor data_in(171) xor data_in(172) xor data_in(173) xor data_in(175) xor data_in(176) xor data_in(180) xor data_in(182) xor data_in(183) xor data_in(188) xor data_in(190) xor data_in(192) xor data_in(194) xor data_in(196) xor data_in(197) xor data_in(199) xor data_in(200) xor data_in(202) xor data_in(204) xor data_in(205) xor data_in(209) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(220) xor data_in(223) xor data_in(224) xor data_in(227) xor data_in(229) xor data_in(238) xor data_in(241) xor data_in(242) xor data_in(244) xor data_in(245) xor data_in(247) xor data_in(252) xor data_in(256) xor data_in(258) xor data_in(260) xor data_in(262) xor data_in(263) xor data_in(265) xor data_in(267) xor data_in(270) xor data_in(271) xor data_in(275) xor data_in(276) xor data_in(277) xor data_in(280) xor data_in(281) xor data_in(283) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(293) xor data_in(295) xor data_in(298) xor data_in(301) xor data_in(303) xor data_in(305) xor data_in(306) xor data_in(309) xor data_in(311) xor data_in(313) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(318) xor data_in(322) xor data_in(323) xor data_in(326) xor data_in(328) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(335) xor data_in(336) xor data_in(338) xor data_in(339) xor data_in(341) xor data_in(342) xor data_in(343) xor data_in(344) xor data_in(347) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(354) xor data_in(356) xor data_in(359) xor data_in(360) xor data_in(362) xor data_in(363) xor data_in(365) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(379) xor data_in(380) xor data_in(381) xor data_in(384) xor data_in(385) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(394) xor data_in(398) xor data_in(399) xor data_in(402) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(420) xor data_in(422) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(429) xor data_in(430) xor data_in(432) xor data_in(433) xor data_in(434) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(444) xor data_in(449) xor data_in(451) xor data_in(452) xor data_in(453) xor data_in(455) xor data_in(456) xor data_in(459) xor data_in(460) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(468) xor data_in(470) xor data_in(471) xor data_in(472) xor data_in(473) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(478) xor data_in(479) xor data_in(480) xor data_in(484) xor data_in(487) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(495) xor data_in(496) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(503) xor data_in(504) xor data_in(507);
    crc_out(3) <= crc_in(2) xor crc_in(5) xor crc_in(6) xor crc_in(9) xor crc_in(10) xor crc_in(14) xor crc_in(17) xor crc_in(18) xor crc_in(22) xor crc_in(23) xor crc_in(24) xor crc_in(27) xor crc_in(33) xor crc_in(35) xor crc_in(37) xor crc_in(39) xor crc_in(42) xor crc_in(50) xor crc_in(51) xor crc_in(54) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(2) xor data_in(5) xor data_in(6) xor data_in(9) xor data_in(10) xor data_in(14) xor data_in(17) xor data_in(18) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(27) xor data_in(33) xor data_in(35) xor data_in(37) xor data_in(39) xor data_in(42) xor data_in(50) xor data_in(51) xor data_in(54) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(65) xor data_in(70) xor data_in(71) xor data_in(74) xor data_in(78) xor data_in(82) xor data_in(84) xor data_in(85) xor data_in(87) xor data_in(89) xor data_in(90) xor data_in(93) xor data_in(95) xor data_in(96) xor data_in(98) xor data_in(103) xor data_in(104) xor data_in(106) xor data_in(107) xor data_in(109) xor data_in(112) xor data_in(113) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(124) xor data_in(126) xor data_in(129) xor data_in(130) xor data_in(131) xor data_in(132) xor data_in(135) xor data_in(137) xor data_in(138) xor data_in(145) xor data_in(146) xor data_in(147) xor data_in(149) xor data_in(151) xor data_in(152) xor data_in(154) xor data_in(156) xor data_in(160) xor data_in(163) xor data_in(165) xor data_in(166) xor data_in(170) xor data_in(172) xor data_in(173) xor data_in(174) xor data_in(176) xor data_in(177) xor data_in(181) xor data_in(183) xor data_in(184) xor data_in(189) xor data_in(191) xor data_in(193) xor data_in(195) xor data_in(197) xor data_in(198) xor data_in(200) xor data_in(201) xor data_in(203) xor data_in(205) xor data_in(206) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(221) xor data_in(224) xor data_in(225) xor data_in(228) xor data_in(230) xor data_in(239) xor data_in(242) xor data_in(243) xor data_in(245) xor data_in(246) xor data_in(248) xor data_in(253) xor data_in(257) xor data_in(259) xor data_in(261) xor data_in(263) xor data_in(264) xor data_in(266) xor data_in(268) xor data_in(271) xor data_in(272) xor data_in(276) xor data_in(277) xor data_in(278) xor data_in(281) xor data_in(282) xor data_in(284) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(294) xor data_in(296) xor data_in(299) xor data_in(302) xor data_in(304) xor data_in(306) xor data_in(307) xor data_in(310) xor data_in(312) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(319) xor data_in(323) xor data_in(324) xor data_in(327) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(340) xor data_in(342) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(348) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(357) xor data_in(360) xor data_in(361) xor data_in(363) xor data_in(364) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(380) xor data_in(381) xor data_in(382) xor data_in(385) xor data_in(386) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(395) xor data_in(399) xor data_in(400) xor data_in(403) xor data_in(406) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(421) xor data_in(423) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(430) xor data_in(431) xor data_in(433) xor data_in(434) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(445) xor data_in(450) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(456) xor data_in(457) xor data_in(460) xor data_in(461) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(469) xor data_in(471) xor data_in(472) xor data_in(473) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(479) xor data_in(480) xor data_in(481) xor data_in(485) xor data_in(488) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(496) xor data_in(497) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(504) xor data_in(505) xor data_in(508);
    crc_out(4) <= crc_in(0) xor crc_in(3) xor crc_in(6) xor crc_in(7) xor crc_in(10) xor crc_in(11) xor crc_in(15) xor crc_in(18) xor crc_in(19) xor crc_in(23) xor crc_in(24) xor crc_in(25) xor crc_in(28) xor crc_in(34) xor crc_in(36) xor crc_in(38) xor crc_in(40) xor crc_in(43) xor crc_in(51) xor crc_in(52) xor crc_in(55) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(3) xor data_in(6) xor data_in(7) xor data_in(10) xor data_in(11) xor data_in(15) xor data_in(18) xor data_in(19) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(28) xor data_in(34) xor data_in(36) xor data_in(38) xor data_in(40) xor data_in(43) xor data_in(51) xor data_in(52) xor data_in(55) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(64) xor data_in(66) xor data_in(71) xor data_in(72) xor data_in(75) xor data_in(79) xor data_in(83) xor data_in(85) xor data_in(86) xor data_in(88) xor data_in(90) xor data_in(91) xor data_in(94) xor data_in(96) xor data_in(97) xor data_in(99) xor data_in(104) xor data_in(105) xor data_in(107) xor data_in(108) xor data_in(110) xor data_in(113) xor data_in(114) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(125) xor data_in(127) xor data_in(130) xor data_in(131) xor data_in(132) xor data_in(133) xor data_in(136) xor data_in(138) xor data_in(139) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(150) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(157) xor data_in(161) xor data_in(164) xor data_in(166) xor data_in(167) xor data_in(171) xor data_in(173) xor data_in(174) xor data_in(175) xor data_in(177) xor data_in(178) xor data_in(182) xor data_in(184) xor data_in(185) xor data_in(190) xor data_in(192) xor data_in(194) xor data_in(196) xor data_in(198) xor data_in(199) xor data_in(201) xor data_in(202) xor data_in(204) xor data_in(206) xor data_in(207) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(222) xor data_in(225) xor data_in(226) xor data_in(229) xor data_in(231) xor data_in(240) xor data_in(243) xor data_in(244) xor data_in(246) xor data_in(247) xor data_in(249) xor data_in(254) xor data_in(258) xor data_in(260) xor data_in(262) xor data_in(264) xor data_in(265) xor data_in(267) xor data_in(269) xor data_in(272) xor data_in(273) xor data_in(277) xor data_in(278) xor data_in(279) xor data_in(282) xor data_in(283) xor data_in(285) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(295) xor data_in(297) xor data_in(300) xor data_in(303) xor data_in(305) xor data_in(307) xor data_in(308) xor data_in(311) xor data_in(313) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(320) xor data_in(324) xor data_in(325) xor data_in(328) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(337) xor data_in(338) xor data_in(340) xor data_in(341) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(349) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(358) xor data_in(361) xor data_in(362) xor data_in(364) xor data_in(365) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(386) xor data_in(387) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(396) xor data_in(400) xor data_in(401) xor data_in(404) xor data_in(407) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(420) xor data_in(422) xor data_in(424) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(431) xor data_in(432) xor data_in(434) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(446) xor data_in(451) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(457) xor data_in(458) xor data_in(461) xor data_in(462) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(470) xor data_in(472) xor data_in(473) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(478) xor data_in(480) xor data_in(481) xor data_in(482) xor data_in(486) xor data_in(489) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(497) xor data_in(498) xor data_in(501) xor data_in(502) xor data_in(503) xor data_in(505) xor data_in(506) xor data_in(509);
    crc_out(5) <= crc_in(0) xor crc_in(1) xor crc_in(4) xor crc_in(7) xor crc_in(8) xor crc_in(11) xor crc_in(12) xor crc_in(16) xor crc_in(19) xor crc_in(20) xor crc_in(24) xor crc_in(25) xor crc_in(26) xor crc_in(29) xor crc_in(35) xor crc_in(37) xor crc_in(39) xor crc_in(41) xor crc_in(44) xor crc_in(52) xor crc_in(53) xor crc_in(56) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(4) xor data_in(7) xor data_in(8) xor data_in(11) xor data_in(12) xor data_in(16) xor data_in(19) xor data_in(20) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(29) xor data_in(35) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(44) xor data_in(52) xor data_in(53) xor data_in(56) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(64) xor data_in(65) xor data_in(67) xor data_in(72) xor data_in(73) xor data_in(76) xor data_in(80) xor data_in(84) xor data_in(86) xor data_in(87) xor data_in(89) xor data_in(91) xor data_in(92) xor data_in(95) xor data_in(97) xor data_in(98) xor data_in(100) xor data_in(105) xor data_in(106) xor data_in(108) xor data_in(109) xor data_in(111) xor data_in(114) xor data_in(115) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(126) xor data_in(128) xor data_in(131) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(137) xor data_in(139) xor data_in(140) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(153) xor data_in(154) xor data_in(156) xor data_in(158) xor data_in(162) xor data_in(165) xor data_in(167) xor data_in(168) xor data_in(172) xor data_in(174) xor data_in(175) xor data_in(176) xor data_in(178) xor data_in(179) xor data_in(183) xor data_in(185) xor data_in(186) xor data_in(191) xor data_in(193) xor data_in(195) xor data_in(197) xor data_in(199) xor data_in(200) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(207) xor data_in(208) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(223) xor data_in(226) xor data_in(227) xor data_in(230) xor data_in(232) xor data_in(241) xor data_in(244) xor data_in(245) xor data_in(247) xor data_in(248) xor data_in(250) xor data_in(255) xor data_in(259) xor data_in(261) xor data_in(263) xor data_in(265) xor data_in(266) xor data_in(268) xor data_in(270) xor data_in(273) xor data_in(274) xor data_in(278) xor data_in(279) xor data_in(280) xor data_in(283) xor data_in(284) xor data_in(286) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(296) xor data_in(298) xor data_in(301) xor data_in(304) xor data_in(306) xor data_in(308) xor data_in(309) xor data_in(312) xor data_in(314) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(321) xor data_in(325) xor data_in(326) xor data_in(329) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(338) xor data_in(339) xor data_in(341) xor data_in(342) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(350) xor data_in(352) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(359) xor data_in(362) xor data_in(363) xor data_in(365) xor data_in(366) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(387) xor data_in(388) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(397) xor data_in(401) xor data_in(402) xor data_in(405) xor data_in(408) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(420) xor data_in(421) xor data_in(423) xor data_in(425) xor data_in(427) xor data_in(428) xor data_in(429) xor data_in(432) xor data_in(433) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(447) xor data_in(452) xor data_in(454) xor data_in(455) xor data_in(456) xor data_in(458) xor data_in(459) xor data_in(462) xor data_in(463) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(471) xor data_in(473) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(481) xor data_in(482) xor data_in(483) xor data_in(487) xor data_in(490) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(498) xor data_in(499) xor data_in(502) xor data_in(503) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(510);
    crc_out(6) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(5) xor crc_in(8) xor crc_in(9) xor crc_in(12) xor crc_in(13) xor crc_in(17) xor crc_in(20) xor crc_in(21) xor crc_in(25) xor crc_in(26) xor crc_in(27) xor crc_in(30) xor crc_in(36) xor crc_in(38) xor crc_in(40) xor crc_in(42) xor crc_in(45) xor crc_in(53) xor crc_in(54) xor crc_in(57) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(5) xor data_in(8) xor data_in(9) xor data_in(12) xor data_in(13) xor data_in(17) xor data_in(20) xor data_in(21) xor data_in(25) xor data_in(26) xor data_in(27) xor data_in(30) xor data_in(36) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(45) xor data_in(53) xor data_in(54) xor data_in(57) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(64) xor data_in(65) xor data_in(66) xor data_in(68) xor data_in(73) xor data_in(74) xor data_in(77) xor data_in(81) xor data_in(85) xor data_in(87) xor data_in(88) xor data_in(90) xor data_in(92) xor data_in(93) xor data_in(96) xor data_in(98) xor data_in(99) xor data_in(101) xor data_in(106) xor data_in(107) xor data_in(109) xor data_in(110) xor data_in(112) xor data_in(115) xor data_in(116) xor data_in(118) xor data_in(119) xor data_in(120) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(127) xor data_in(129) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(138) xor data_in(140) xor data_in(141) xor data_in(148) xor data_in(149) xor data_in(150) xor data_in(152) xor data_in(154) xor data_in(155) xor data_in(157) xor data_in(159) xor data_in(163) xor data_in(166) xor data_in(168) xor data_in(169) xor data_in(173) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(179) xor data_in(180) xor data_in(184) xor data_in(186) xor data_in(187) xor data_in(192) xor data_in(194) xor data_in(196) xor data_in(198) xor data_in(200) xor data_in(201) xor data_in(203) xor data_in(204) xor data_in(206) xor data_in(208) xor data_in(209) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(224) xor data_in(227) xor data_in(228) xor data_in(231) xor data_in(233) xor data_in(242) xor data_in(245) xor data_in(246) xor data_in(248) xor data_in(249) xor data_in(251) xor data_in(256) xor data_in(260) xor data_in(262) xor data_in(264) xor data_in(266) xor data_in(267) xor data_in(269) xor data_in(271) xor data_in(274) xor data_in(275) xor data_in(279) xor data_in(280) xor data_in(281) xor data_in(284) xor data_in(285) xor data_in(287) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(295) xor data_in(297) xor data_in(299) xor data_in(302) xor data_in(305) xor data_in(307) xor data_in(309) xor data_in(310) xor data_in(313) xor data_in(315) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(322) xor data_in(326) xor data_in(327) xor data_in(330) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(339) xor data_in(340) xor data_in(342) xor data_in(343) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(351) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(360) xor data_in(363) xor data_in(364) xor data_in(366) xor data_in(367) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(383) xor data_in(384) xor data_in(385) xor data_in(388) xor data_in(389) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(398) xor data_in(402) xor data_in(403) xor data_in(406) xor data_in(409) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(420) xor data_in(421) xor data_in(422) xor data_in(424) xor data_in(426) xor data_in(428) xor data_in(429) xor data_in(430) xor data_in(433) xor data_in(434) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(448) xor data_in(453) xor data_in(455) xor data_in(456) xor data_in(457) xor data_in(459) xor data_in(460) xor data_in(463) xor data_in(464) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(472) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(480) xor data_in(482) xor data_in(483) xor data_in(484) xor data_in(488) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(499) xor data_in(500) xor data_in(503) xor data_in(504) xor data_in(505) xor data_in(507) xor data_in(508) xor data_in(511);
    crc_out(7) <= crc_in(0) xor crc_in(1) xor crc_in(3) xor crc_in(5) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(12) xor crc_in(15) xor crc_in(18) xor crc_in(24) xor crc_in(26) xor crc_in(27) xor crc_in(28) xor crc_in(31) xor crc_in(32) xor crc_in(36) xor crc_in(37) xor crc_in(39) xor crc_in(45) xor crc_in(46) xor crc_in(47) xor crc_in(50) xor crc_in(52) xor crc_in(53) xor crc_in(59) xor crc_in(61) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(12) xor data_in(15) xor data_in(18) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(31) xor data_in(32) xor data_in(36) xor data_in(37) xor data_in(39) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(50) xor data_in(52) xor data_in(53) xor data_in(59) xor data_in(61) xor data_in(63) xor data_in(64) xor data_in(65) xor data_in(66) xor data_in(67) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(79) xor data_in(80) xor data_in(83) xor data_in(85) xor data_in(87) xor data_in(88) xor data_in(89) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(97) xor data_in(99) xor data_in(100) xor data_in(103) xor data_in(104) xor data_in(107) xor data_in(114) xor data_in(116) xor data_in(117) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(125) xor data_in(128) xor data_in(129) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(137) xor data_in(138) xor data_in(140) xor data_in(143) xor data_in(146) xor data_in(149) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(157) xor data_in(165) xor data_in(166) xor data_in(168) xor data_in(169) xor data_in(171) xor data_in(174) xor data_in(175) xor data_in(179) xor data_in(180) xor data_in(182) xor data_in(184) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(190) xor data_in(193) xor data_in(194) xor data_in(195) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(206) xor data_in(208) xor data_in(209) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(215) xor data_in(217) xor data_in(223) xor data_in(224) xor data_in(226) xor data_in(230) xor data_in(231) xor data_in(233) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(239) xor data_in(242) xor data_in(243) xor data_in(245) xor data_in(246) xor data_in(247) xor data_in(249) xor data_in(250) xor data_in(254) xor data_in(257) xor data_in(258) xor data_in(261) xor data_in(262) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(278) xor data_in(280) xor data_in(282) xor data_in(285) xor data_in(286) xor data_in(287) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(296) xor data_in(297) xor data_in(299) xor data_in(302) xor data_in(304) xor data_in(306) xor data_in(308) xor data_in(309) xor data_in(310) xor data_in(311) xor data_in(313) xor data_in(316) xor data_in(319) xor data_in(321) xor data_in(325) xor data_in(326) xor data_in(328) xor data_in(330) xor data_in(332) xor data_in(335) xor data_in(336) xor data_in(338) xor data_in(339) xor data_in(341) xor data_in(345) xor data_in(347) xor data_in(353) xor data_in(354) xor data_in(359) xor data_in(361) xor data_in(362) xor data_in(363) xor data_in(365) xor data_in(370) xor data_in(371) xor data_in(374) xor data_in(375) xor data_in(377) xor data_in(378) xor data_in(382) xor data_in(384) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(394) xor data_in(396) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(414) xor data_in(415) xor data_in(418) xor data_in(422) xor data_in(424) xor data_in(425) xor data_in(427) xor data_in(437) xor data_in(440) xor data_in(441) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(452) xor data_in(453) xor data_in(456) xor data_in(457) xor data_in(458) xor data_in(459) xor data_in(462) xor data_in(463) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(469) xor data_in(473) xor data_in(474) xor data_in(476) xor data_in(479) xor data_in(480) xor data_in(481) xor data_in(483) xor data_in(485) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(498) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(503) xor data_in(509) xor data_in(510);
    crc_out(8) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(4) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(10) xor crc_in(13) xor crc_in(16) xor crc_in(19) xor crc_in(25) xor crc_in(27) xor crc_in(28) xor crc_in(29) xor crc_in(32) xor crc_in(33) xor crc_in(37) xor crc_in(38) xor crc_in(40) xor crc_in(46) xor crc_in(47) xor crc_in(48) xor crc_in(51) xor crc_in(53) xor crc_in(54) xor crc_in(60) xor crc_in(62) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(13) xor data_in(16) xor data_in(19) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(32) xor data_in(33) xor data_in(37) xor data_in(38) xor data_in(40) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(53) xor data_in(54) xor data_in(60) xor data_in(62) xor data_in(64) xor data_in(65) xor data_in(66) xor data_in(67) xor data_in(68) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(76) xor data_in(77) xor data_in(78) xor data_in(80) xor data_in(81) xor data_in(84) xor data_in(86) xor data_in(88) xor data_in(89) xor data_in(90) xor data_in(92) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(98) xor data_in(100) xor data_in(101) xor data_in(104) xor data_in(105) xor data_in(108) xor data_in(115) xor data_in(117) xor data_in(118) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(126) xor data_in(129) xor data_in(130) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(136) xor data_in(138) xor data_in(139) xor data_in(141) xor data_in(144) xor data_in(147) xor data_in(150) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(158) xor data_in(166) xor data_in(167) xor data_in(169) xor data_in(170) xor data_in(172) xor data_in(175) xor data_in(176) xor data_in(180) xor data_in(181) xor data_in(183) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(191) xor data_in(194) xor data_in(195) xor data_in(196) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(207) xor data_in(209) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(216) xor data_in(218) xor data_in(224) xor data_in(225) xor data_in(227) xor data_in(231) xor data_in(232) xor data_in(234) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(240) xor data_in(243) xor data_in(244) xor data_in(246) xor data_in(247) xor data_in(248) xor data_in(250) xor data_in(251) xor data_in(255) xor data_in(258) xor data_in(259) xor data_in(262) xor data_in(263) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(279) xor data_in(281) xor data_in(283) xor data_in(286) xor data_in(287) xor data_in(288) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(295) xor data_in(297) xor data_in(298) xor data_in(300) xor data_in(303) xor data_in(305) xor data_in(307) xor data_in(309) xor data_in(310) xor data_in(311) xor data_in(312) xor data_in(314) xor data_in(317) xor data_in(320) xor data_in(322) xor data_in(326) xor data_in(327) xor data_in(329) xor data_in(331) xor data_in(333) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(340) xor data_in(342) xor data_in(346) xor data_in(348) xor data_in(354) xor data_in(355) xor data_in(360) xor data_in(362) xor data_in(363) xor data_in(364) xor data_in(366) xor data_in(371) xor data_in(372) xor data_in(375) xor data_in(376) xor data_in(378) xor data_in(379) xor data_in(383) xor data_in(385) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(395) xor data_in(397) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(415) xor data_in(416) xor data_in(419) xor data_in(423) xor data_in(425) xor data_in(426) xor data_in(428) xor data_in(438) xor data_in(441) xor data_in(442) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(453) xor data_in(454) xor data_in(457) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(463) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(470) xor data_in(474) xor data_in(475) xor data_in(477) xor data_in(480) xor data_in(481) xor data_in(482) xor data_in(484) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(490) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(504) xor data_in(510) xor data_in(511);
    crc_out(9) <= crc_in(1) xor crc_in(3) xor crc_in(9) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(15) xor crc_in(17) xor crc_in(20) xor crc_in(21) xor crc_in(22) xor crc_in(24) xor crc_in(26) xor crc_in(28) xor crc_in(29) xor crc_in(30) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(36) xor crc_in(38) xor crc_in(39) xor crc_in(43) xor crc_in(45) xor crc_in(48) xor crc_in(49) xor crc_in(50) xor crc_in(53) xor crc_in(58) xor crc_in(59) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(1) xor data_in(3) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(17) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(24) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(36) xor data_in(38) xor data_in(39) xor data_in(43) xor data_in(45) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(53) xor data_in(58) xor data_in(59) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(65) xor data_in(66) xor data_in(67) xor data_in(68) xor data_in(70) xor data_in(71) xor data_in(73) xor data_in(76) xor data_in(80) xor data_in(81) xor data_in(83) xor data_in(86) xor data_in(89) xor data_in(90) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(94) xor data_in(96) xor data_in(97) xor data_in(99) xor data_in(101) xor data_in(103) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(111) xor data_in(113) xor data_in(114) xor data_in(116) xor data_in(118) xor data_in(120) xor data_in(122) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(129) xor data_in(131) xor data_in(132) xor data_in(134) xor data_in(135) xor data_in(138) xor data_in(141) xor data_in(143) xor data_in(145) xor data_in(146) xor data_in(148) xor data_in(150) xor data_in(152) xor data_in(157) xor data_in(158) xor data_in(159) xor data_in(160) xor data_in(164) xor data_in(165) xor data_in(166) xor data_in(173) xor data_in(175) xor data_in(178) xor data_in(179) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(192) xor data_in(194) xor data_in(195) xor data_in(196) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(210) xor data_in(213) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(223) xor data_in(224) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(234) xor data_in(236) xor data_in(238) xor data_in(241) xor data_in(242) xor data_in(244) xor data_in(247) xor data_in(248) xor data_in(249) xor data_in(251) xor data_in(254) xor data_in(256) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(262) xor data_in(269) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(275) xor data_in(276) xor data_in(278) xor data_in(280) xor data_in(281) xor data_in(282) xor data_in(284) xor data_in(289) xor data_in(291) xor data_in(293) xor data_in(294) xor data_in(296) xor data_in(297) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(306) xor data_in(308) xor data_in(309) xor data_in(310) xor data_in(311) xor data_in(312) xor data_in(314) xor data_in(315) xor data_in(320) xor data_in(321) xor data_in(325) xor data_in(326) xor data_in(328) xor data_in(331) xor data_in(333) xor data_in(337) xor data_in(339) xor data_in(341) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(352) xor data_in(353) xor data_in(357) xor data_in(358) xor data_in(361) xor data_in(362) xor data_in(365) xor data_in(368) xor data_in(376) xor data_in(377) xor data_in(382) xor data_in(384) xor data_in(385) xor data_in(386) xor data_in(387) xor data_in(389) xor data_in(390) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(401) xor data_in(402) xor data_in(406) xor data_in(407) xor data_in(408) xor data_in(410) xor data_in(411) xor data_in(413) xor data_in(419) xor data_in(421) xor data_in(423) xor data_in(426) xor data_in(427) xor data_in(430) xor data_in(431) xor data_in(434) xor data_in(435) xor data_in(438) xor data_in(443) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(452) xor data_in(453) xor data_in(455) xor data_in(458) xor data_in(462) xor data_in(463) xor data_in(464) xor data_in(465) xor data_in(467) xor data_in(468) xor data_in(470) xor data_in(474) xor data_in(476) xor data_in(477) xor data_in(481) xor data_in(482) xor data_in(483) xor data_in(484) xor data_in(485) xor data_in(486) xor data_in(489) xor data_in(490) xor data_in(494) xor data_in(495) xor data_in(497) xor data_in(498) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(504) xor data_in(506) xor data_in(508) xor data_in(510) xor data_in(511);
    crc_out(10) <= crc_in(4) xor crc_in(5) xor crc_in(7) xor crc_in(8) xor crc_in(15) xor crc_in(16) xor crc_in(18) xor crc_in(23) xor crc_in(24) xor crc_in(25) xor crc_in(27) xor crc_in(29) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(37) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(47) xor crc_in(49) xor crc_in(51) xor crc_in(52) xor crc_in(53) xor crc_in(55) xor crc_in(58) xor crc_in(60) xor crc_in(63) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(49) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(58) xor data_in(60) xor data_in(63) xor data_in(64) xor data_in(66) xor data_in(67) xor data_in(68) xor data_in(70) xor data_in(76) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(90) xor data_in(91) xor data_in(93) xor data_in(94) xor data_in(97) xor data_in(98) xor data_in(100) xor data_in(103) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(112) xor data_in(113) xor data_in(115) xor data_in(117) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(124) xor data_in(127) xor data_in(128) xor data_in(129) xor data_in(133) xor data_in(135) xor data_in(137) xor data_in(138) xor data_in(140) xor data_in(141) xor data_in(143) xor data_in(144) xor data_in(147) xor data_in(149) xor data_in(150) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(159) xor data_in(161) xor data_in(164) xor data_in(168) xor data_in(170) xor data_in(171) xor data_in(174) xor data_in(175) xor data_in(177) xor data_in(178) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(184) xor data_in(186) xor data_in(188) xor data_in(189) xor data_in(193) xor data_in(194) xor data_in(195) xor data_in(196) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(212) xor data_in(216) xor data_in(217) xor data_in(219) xor data_in(220) xor data_in(223) xor data_in(226) xor data_in(228) xor data_in(229) xor data_in(233) xor data_in(234) xor data_in(236) xor data_in(243) xor data_in(248) xor data_in(249) xor data_in(250) xor data_in(254) xor data_in(255) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(262) xor data_in(264) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(273) xor data_in(277) xor data_in(278) xor data_in(279) xor data_in(282) xor data_in(283) xor data_in(285) xor data_in(287) xor data_in(288) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(294) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(307) xor data_in(310) xor data_in(311) xor data_in(312) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(318) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(325) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(333) xor data_in(339) xor data_in(342) xor data_in(343) xor data_in(344) xor data_in(347) xor data_in(352) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(359) xor data_in(364) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(372) xor data_in(373) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(380) xor data_in(382) xor data_in(383) xor data_in(386) xor data_in(390) xor data_in(392) xor data_in(393) xor data_in(396) xor data_in(400) xor data_in(402) xor data_in(403) xor data_in(405) xor data_in(407) xor data_in(411) xor data_in(413) xor data_in(414) xor data_in(416) xor data_in(417) xor data_in(419) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(427) xor data_in(428) xor data_in(429) xor data_in(430) xor data_in(432) xor data_in(434) xor data_in(436) xor data_in(438) xor data_in(442) xor data_in(444) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(452) xor data_in(456) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(464) xor data_in(465) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(474) xor data_in(482) xor data_in(483) xor data_in(485) xor data_in(488) xor data_in(490) xor data_in(493) xor data_in(495) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(509) xor data_in(510) xor data_in(511);
    crc_out(11) <= crc_in(2) xor crc_in(6) xor crc_in(7) xor crc_in(9) xor crc_in(10) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(17) xor crc_in(19) xor crc_in(21) xor crc_in(22) xor crc_in(25) xor crc_in(26) xor crc_in(28) xor crc_in(30) xor crc_in(31) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(37) xor crc_in(38) xor crc_in(40) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(46) xor crc_in(48) xor crc_in(55) xor crc_in(56) xor crc_in(58) xor crc_in(61) xor crc_in(62) xor data_in(2) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(37) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(48) xor data_in(55) xor data_in(56) xor data_in(58) xor data_in(61) xor data_in(62) xor data_in(64) xor data_in(65) xor data_in(67) xor data_in(68) xor data_in(70) xor data_in(72) xor data_in(74) xor data_in(76) xor data_in(78) xor data_in(81) xor data_in(83) xor data_in(84) xor data_in(91) xor data_in(94) xor data_in(98) xor data_in(99) xor data_in(101) xor data_in(102) xor data_in(103) xor data_in(106) xor data_in(107) xor data_in(109) xor data_in(111) xor data_in(116) xor data_in(118) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(124) xor data_in(125) xor data_in(126) xor data_in(128) xor data_in(132) xor data_in(134) xor data_in(137) xor data_in(140) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(148) xor data_in(152) xor data_in(153) xor data_in(162) xor data_in(164) xor data_in(166) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(170) xor data_in(172) xor data_in(177) xor data_in(183) xor data_in(184) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(189) xor data_in(195) xor data_in(196) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(207) xor data_in(208) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(216) xor data_in(217) xor data_in(220) xor data_in(221) xor data_in(223) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(236) xor data_in(239) xor data_in(242) xor data_in(244) xor data_in(245) xor data_in(249) xor data_in(250) xor data_in(251) xor data_in(252) xor data_in(254) xor data_in(255) xor data_in(256) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(274) xor data_in(275) xor data_in(276) xor data_in(279) xor data_in(280) xor data_in(281) xor data_in(283) xor data_in(284) xor data_in(286) xor data_in(287) xor data_in(289) xor data_in(292) xor data_in(293) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(301) xor data_in(303) xor data_in(304) xor data_in(308) xor data_in(309) xor data_in(311) xor data_in(312) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(324) xor data_in(325) xor data_in(327) xor data_in(333) xor data_in(338) xor data_in(339) xor data_in(346) xor data_in(349) xor data_in(352) xor data_in(360) xor data_in(362) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(369) xor data_in(370) xor data_in(372) xor data_in(374) xor data_in(378) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(385) xor data_in(388) xor data_in(392) xor data_in(394) xor data_in(395) xor data_in(398) xor data_in(400) xor data_in(401) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(409) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(418) xor data_in(419) xor data_in(421) xor data_in(422) xor data_in(428) xor data_in(433) xor data_in(434) xor data_in(437) xor data_in(438) xor data_in(442) xor data_in(443) xor data_in(445) xor data_in(447) xor data_in(448) xor data_in(452) xor data_in(454) xor data_in(457) xor data_in(459) xor data_in(460) xor data_in(465) xor data_in(469) xor data_in(474) xor data_in(477) xor data_in(478) xor data_in(483) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(493) xor data_in(494) xor data_in(498) xor data_in(499) xor data_in(501) xor data_in(502) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(509) xor data_in(511);
    crc_out(12) <= crc_in(2) xor crc_in(3) xor crc_in(5) xor crc_in(11) xor crc_in(12) xor crc_in(16) xor crc_in(17) xor crc_in(18) xor crc_in(20) xor crc_in(21) xor crc_in(23) xor crc_in(24) xor crc_in(26) xor crc_in(27) xor crc_in(29) xor crc_in(31) xor crc_in(34) xor crc_in(35) xor crc_in(38) xor crc_in(39) xor crc_in(44) xor crc_in(49) xor crc_in(50) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(63) xor data_in(2) xor data_in(3) xor data_in(5) xor data_in(11) xor data_in(12) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(29) xor data_in(31) xor data_in(34) xor data_in(35) xor data_in(38) xor data_in(39) xor data_in(44) xor data_in(49) xor data_in(50) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(63) xor data_in(65) xor data_in(66) xor data_in(68) xor data_in(70) xor data_in(72) xor data_in(73) xor data_in(74) xor data_in(75) xor data_in(76) xor data_in(78) xor data_in(80) xor data_in(83) xor data_in(84) xor data_in(86) xor data_in(87) xor data_in(99) xor data_in(100) xor data_in(107) xor data_in(111) xor data_in(112) xor data_in(113) xor data_in(114) xor data_in(117) xor data_in(121) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(127) xor data_in(130) xor data_in(132) xor data_in(133) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(139) xor data_in(140) xor data_in(142) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(147) xor data_in(149) xor data_in(150) xor data_in(151) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(158) xor data_in(160) xor data_in(163) xor data_in(164) xor data_in(166) xor data_in(169) xor data_in(173) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(179) xor data_in(181) xor data_in(182) xor data_in(185) xor data_in(187) xor data_in(188) xor data_in(194) xor data_in(196) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(207) xor data_in(209) xor data_in(211) xor data_in(213) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(221) xor data_in(222) xor data_in(223) xor data_in(225) xor data_in(227) xor data_in(230) xor data_in(231) xor data_in(235) xor data_in(236) xor data_in(239) xor data_in(240) xor data_in(242) xor data_in(243) xor data_in(246) xor data_in(250) xor data_in(251) xor data_in(253) xor data_in(254) xor data_in(255) xor data_in(256) xor data_in(257) xor data_in(258) xor data_in(260) xor data_in(261) xor data_in(263) xor data_in(264) xor data_in(265) xor data_in(268) xor data_in(269) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(277) xor data_in(278) xor data_in(280) xor data_in(282) xor data_in(284) xor data_in(285) xor data_in(290) xor data_in(291) xor data_in(293) xor data_in(294) xor data_in(295) xor data_in(297) xor data_in(303) xor data_in(305) xor data_in(310) xor data_in(312) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(319) xor data_in(321) xor data_in(322) xor data_in(327) xor data_in(328) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(338) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(352) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(361) xor data_in(362) xor data_in(365) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(375) xor data_in(380) xor data_in(383) xor data_in(384) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(391) xor data_in(392) xor data_in(396) xor data_in(397) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(402) xor data_in(404) xor data_in(406) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(421) xor data_in(422) xor data_in(424) xor data_in(430) xor data_in(431) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(446) xor data_in(448) xor data_in(452) xor data_in(454) xor data_in(455) xor data_in(458) xor data_in(459) xor data_in(462) xor data_in(463) xor data_in(471) xor data_in(474) xor data_in(477) xor data_in(479) xor data_in(486) xor data_in(487) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(498) xor data_in(500) xor data_in(502) xor data_in(504) xor data_in(506) xor data_in(507);
    crc_out(13) <= crc_in(3) xor crc_in(4) xor crc_in(6) xor crc_in(12) xor crc_in(13) xor crc_in(17) xor crc_in(18) xor crc_in(19) xor crc_in(21) xor crc_in(22) xor crc_in(24) xor crc_in(25) xor crc_in(27) xor crc_in(28) xor crc_in(30) xor crc_in(32) xor crc_in(35) xor crc_in(36) xor crc_in(39) xor crc_in(40) xor crc_in(45) xor crc_in(50) xor crc_in(51) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor data_in(3) xor data_in(4) xor data_in(6) xor data_in(12) xor data_in(13) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(32) xor data_in(35) xor data_in(36) xor data_in(39) xor data_in(40) xor data_in(45) xor data_in(50) xor data_in(51) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(64) xor data_in(66) xor data_in(67) xor data_in(69) xor data_in(71) xor data_in(73) xor data_in(74) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(79) xor data_in(81) xor data_in(84) xor data_in(85) xor data_in(87) xor data_in(88) xor data_in(100) xor data_in(101) xor data_in(108) xor data_in(112) xor data_in(113) xor data_in(114) xor data_in(115) xor data_in(118) xor data_in(122) xor data_in(124) xor data_in(125) xor data_in(126) xor data_in(128) xor data_in(131) xor data_in(133) xor data_in(134) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(140) xor data_in(141) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(148) xor data_in(150) xor data_in(151) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(156) xor data_in(157) xor data_in(158) xor data_in(159) xor data_in(161) xor data_in(164) xor data_in(165) xor data_in(167) xor data_in(170) xor data_in(174) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(180) xor data_in(182) xor data_in(183) xor data_in(186) xor data_in(188) xor data_in(189) xor data_in(195) xor data_in(197) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(204) xor data_in(206) xor data_in(208) xor data_in(210) xor data_in(212) xor data_in(214) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(222) xor data_in(223) xor data_in(224) xor data_in(226) xor data_in(228) xor data_in(231) xor data_in(232) xor data_in(236) xor data_in(237) xor data_in(240) xor data_in(241) xor data_in(243) xor data_in(244) xor data_in(247) xor data_in(251) xor data_in(252) xor data_in(254) xor data_in(255) xor data_in(256) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(261) xor data_in(262) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(273) xor data_in(275) xor data_in(278) xor data_in(279) xor data_in(281) xor data_in(283) xor data_in(285) xor data_in(286) xor data_in(291) xor data_in(292) xor data_in(294) xor data_in(295) xor data_in(296) xor data_in(298) xor data_in(304) xor data_in(306) xor data_in(311) xor data_in(313) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(320) xor data_in(322) xor data_in(323) xor data_in(328) xor data_in(329) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(339) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(353) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(362) xor data_in(363) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(376) xor data_in(381) xor data_in(384) xor data_in(385) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(392) xor data_in(393) xor data_in(397) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(402) xor data_in(403) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(422) xor data_in(423) xor data_in(425) xor data_in(431) xor data_in(432) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(447) xor data_in(449) xor data_in(453) xor data_in(455) xor data_in(456) xor data_in(459) xor data_in(460) xor data_in(463) xor data_in(464) xor data_in(472) xor data_in(475) xor data_in(478) xor data_in(480) xor data_in(487) xor data_in(488) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(497) xor data_in(499) xor data_in(501) xor data_in(503) xor data_in(505) xor data_in(507) xor data_in(508);
    crc_out(14) <= crc_in(0) xor crc_in(4) xor crc_in(5) xor crc_in(7) xor crc_in(13) xor crc_in(14) xor crc_in(18) xor crc_in(19) xor crc_in(20) xor crc_in(22) xor crc_in(23) xor crc_in(25) xor crc_in(26) xor crc_in(28) xor crc_in(29) xor crc_in(31) xor crc_in(33) xor crc_in(36) xor crc_in(37) xor crc_in(40) xor crc_in(41) xor crc_in(46) xor crc_in(51) xor crc_in(52) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor data_in(0) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(13) xor data_in(14) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(33) xor data_in(36) xor data_in(37) xor data_in(40) xor data_in(41) xor data_in(46) xor data_in(51) xor data_in(52) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(65) xor data_in(67) xor data_in(68) xor data_in(70) xor data_in(72) xor data_in(74) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(78) xor data_in(80) xor data_in(82) xor data_in(85) xor data_in(86) xor data_in(88) xor data_in(89) xor data_in(101) xor data_in(102) xor data_in(109) xor data_in(113) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(119) xor data_in(123) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(129) xor data_in(132) xor data_in(134) xor data_in(135) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(141) xor data_in(142) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(147) xor data_in(149) xor data_in(151) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(157) xor data_in(158) xor data_in(159) xor data_in(160) xor data_in(162) xor data_in(165) xor data_in(166) xor data_in(168) xor data_in(171) xor data_in(175) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(181) xor data_in(183) xor data_in(184) xor data_in(187) xor data_in(189) xor data_in(190) xor data_in(196) xor data_in(198) xor data_in(202) xor data_in(203) xor data_in(204) xor data_in(205) xor data_in(207) xor data_in(209) xor data_in(211) xor data_in(213) xor data_in(215) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(223) xor data_in(224) xor data_in(225) xor data_in(227) xor data_in(229) xor data_in(232) xor data_in(233) xor data_in(237) xor data_in(238) xor data_in(241) xor data_in(242) xor data_in(244) xor data_in(245) xor data_in(248) xor data_in(252) xor data_in(253) xor data_in(255) xor data_in(256) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(262) xor data_in(263) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(274) xor data_in(276) xor data_in(279) xor data_in(280) xor data_in(282) xor data_in(284) xor data_in(286) xor data_in(287) xor data_in(292) xor data_in(293) xor data_in(295) xor data_in(296) xor data_in(297) xor data_in(299) xor data_in(305) xor data_in(307) xor data_in(312) xor data_in(314) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(321) xor data_in(323) xor data_in(324) xor data_in(329) xor data_in(330) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(340) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(354) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(363) xor data_in(364) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(377) xor data_in(382) xor data_in(385) xor data_in(386) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(393) xor data_in(394) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(402) xor data_in(403) xor data_in(404) xor data_in(406) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(423) xor data_in(424) xor data_in(426) xor data_in(432) xor data_in(433) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(448) xor data_in(450) xor data_in(454) xor data_in(456) xor data_in(457) xor data_in(460) xor data_in(461) xor data_in(464) xor data_in(465) xor data_in(473) xor data_in(476) xor data_in(479) xor data_in(481) xor data_in(488) xor data_in(489) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(495) xor data_in(496) xor data_in(497) xor data_in(498) xor data_in(500) xor data_in(502) xor data_in(504) xor data_in(506) xor data_in(508) xor data_in(509);
    crc_out(15) <= crc_in(1) xor crc_in(5) xor crc_in(6) xor crc_in(8) xor crc_in(14) xor crc_in(15) xor crc_in(19) xor crc_in(20) xor crc_in(21) xor crc_in(23) xor crc_in(24) xor crc_in(26) xor crc_in(27) xor crc_in(29) xor crc_in(30) xor crc_in(32) xor crc_in(34) xor crc_in(37) xor crc_in(38) xor crc_in(41) xor crc_in(42) xor crc_in(47) xor crc_in(52) xor crc_in(53) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor data_in(1) xor data_in(5) xor data_in(6) xor data_in(8) xor data_in(14) xor data_in(15) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(34) xor data_in(37) xor data_in(38) xor data_in(41) xor data_in(42) xor data_in(47) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(66) xor data_in(68) xor data_in(69) xor data_in(71) xor data_in(73) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(81) xor data_in(83) xor data_in(86) xor data_in(87) xor data_in(89) xor data_in(90) xor data_in(102) xor data_in(103) xor data_in(110) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(120) xor data_in(124) xor data_in(126) xor data_in(127) xor data_in(128) xor data_in(130) xor data_in(133) xor data_in(135) xor data_in(136) xor data_in(138) xor data_in(139) xor data_in(140) xor data_in(142) xor data_in(143) xor data_in(145) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(150) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(156) xor data_in(158) xor data_in(159) xor data_in(160) xor data_in(161) xor data_in(163) xor data_in(166) xor data_in(167) xor data_in(169) xor data_in(172) xor data_in(176) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(182) xor data_in(184) xor data_in(185) xor data_in(188) xor data_in(190) xor data_in(191) xor data_in(197) xor data_in(199) xor data_in(203) xor data_in(204) xor data_in(205) xor data_in(206) xor data_in(208) xor data_in(210) xor data_in(212) xor data_in(214) xor data_in(216) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(224) xor data_in(225) xor data_in(226) xor data_in(228) xor data_in(230) xor data_in(233) xor data_in(234) xor data_in(238) xor data_in(239) xor data_in(242) xor data_in(243) xor data_in(245) xor data_in(246) xor data_in(249) xor data_in(253) xor data_in(254) xor data_in(256) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(263) xor data_in(264) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(275) xor data_in(277) xor data_in(280) xor data_in(281) xor data_in(283) xor data_in(285) xor data_in(287) xor data_in(288) xor data_in(293) xor data_in(294) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(300) xor data_in(306) xor data_in(308) xor data_in(313) xor data_in(315) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(322) xor data_in(324) xor data_in(325) xor data_in(330) xor data_in(331) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(336) xor data_in(341) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(355) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(364) xor data_in(365) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(378) xor data_in(383) xor data_in(386) xor data_in(387) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(394) xor data_in(395) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(402) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(407) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(424) xor data_in(425) xor data_in(427) xor data_in(433) xor data_in(434) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(449) xor data_in(451) xor data_in(455) xor data_in(457) xor data_in(458) xor data_in(461) xor data_in(462) xor data_in(465) xor data_in(466) xor data_in(474) xor data_in(477) xor data_in(480) xor data_in(482) xor data_in(489) xor data_in(490) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(496) xor data_in(497) xor data_in(498) xor data_in(499) xor data_in(501) xor data_in(503) xor data_in(505) xor data_in(507) xor data_in(509) xor data_in(510);
    crc_out(16) <= crc_in(2) xor crc_in(6) xor crc_in(7) xor crc_in(9) xor crc_in(15) xor crc_in(16) xor crc_in(20) xor crc_in(21) xor crc_in(22) xor crc_in(24) xor crc_in(25) xor crc_in(27) xor crc_in(28) xor crc_in(30) xor crc_in(31) xor crc_in(33) xor crc_in(35) xor crc_in(38) xor crc_in(39) xor crc_in(42) xor crc_in(43) xor crc_in(48) xor crc_in(53) xor crc_in(54) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor data_in(2) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(15) xor data_in(16) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(33) xor data_in(35) xor data_in(38) xor data_in(39) xor data_in(42) xor data_in(43) xor data_in(48) xor data_in(53) xor data_in(54) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(67) xor data_in(69) xor data_in(70) xor data_in(72) xor data_in(74) xor data_in(76) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(82) xor data_in(84) xor data_in(87) xor data_in(88) xor data_in(90) xor data_in(91) xor data_in(103) xor data_in(104) xor data_in(111) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(121) xor data_in(125) xor data_in(127) xor data_in(128) xor data_in(129) xor data_in(131) xor data_in(134) xor data_in(136) xor data_in(137) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(143) xor data_in(144) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(159) xor data_in(160) xor data_in(161) xor data_in(162) xor data_in(164) xor data_in(167) xor data_in(168) xor data_in(170) xor data_in(173) xor data_in(177) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(183) xor data_in(185) xor data_in(186) xor data_in(189) xor data_in(191) xor data_in(192) xor data_in(198) xor data_in(200) xor data_in(204) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(209) xor data_in(211) xor data_in(213) xor data_in(215) xor data_in(217) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(229) xor data_in(231) xor data_in(234) xor data_in(235) xor data_in(239) xor data_in(240) xor data_in(243) xor data_in(244) xor data_in(246) xor data_in(247) xor data_in(250) xor data_in(254) xor data_in(255) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(262) xor data_in(264) xor data_in(265) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(272) xor data_in(273) xor data_in(275) xor data_in(276) xor data_in(278) xor data_in(281) xor data_in(282) xor data_in(284) xor data_in(286) xor data_in(288) xor data_in(289) xor data_in(294) xor data_in(295) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(301) xor data_in(307) xor data_in(309) xor data_in(314) xor data_in(316) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(321) xor data_in(323) xor data_in(325) xor data_in(326) xor data_in(331) xor data_in(332) xor data_in(334) xor data_in(335) xor data_in(336) xor data_in(337) xor data_in(342) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(354) xor data_in(356) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(362) xor data_in(365) xor data_in(366) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(379) xor data_in(384) xor data_in(387) xor data_in(388) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(395) xor data_in(396) xor data_in(400) xor data_in(401) xor data_in(402) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(408) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(425) xor data_in(426) xor data_in(428) xor data_in(434) xor data_in(435) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(450) xor data_in(452) xor data_in(456) xor data_in(458) xor data_in(459) xor data_in(462) xor data_in(463) xor data_in(466) xor data_in(467) xor data_in(475) xor data_in(478) xor data_in(481) xor data_in(483) xor data_in(490) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(497) xor data_in(498) xor data_in(499) xor data_in(500) xor data_in(502) xor data_in(504) xor data_in(506) xor data_in(508) xor data_in(510) xor data_in(511);
    crc_out(17) <= crc_in(2) xor crc_in(3) xor crc_in(5) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(17) xor crc_in(23) xor crc_in(24) xor crc_in(25) xor crc_in(26) xor crc_in(28) xor crc_in(29) xor crc_in(31) xor crc_in(34) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(44) xor crc_in(45) xor crc_in(47) xor crc_in(49) xor crc_in(50) xor crc_in(52) xor crc_in(53) xor crc_in(57) xor crc_in(60) xor crc_in(61) xor crc_in(63) xor data_in(2) xor data_in(3) xor data_in(5) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(34) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(49) xor data_in(50) xor data_in(52) xor data_in(53) xor data_in(57) xor data_in(60) xor data_in(61) xor data_in(63) xor data_in(68) xor data_in(69) xor data_in(72) xor data_in(73) xor data_in(74) xor data_in(75) xor data_in(76) xor data_in(81) xor data_in(82) xor data_in(86) xor data_in(87) xor data_in(88) xor data_in(89) xor data_in(91) xor data_in(95) xor data_in(102) xor data_in(103) xor data_in(105) xor data_in(108) xor data_in(110) xor data_in(111) xor data_in(112) xor data_in(113) xor data_in(114) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(120) xor data_in(123) xor data_in(124) xor data_in(128) xor data_in(135) xor data_in(136) xor data_in(139) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(161) xor data_in(162) xor data_in(163) xor data_in(164) xor data_in(166) xor data_in(167) xor data_in(169) xor data_in(170) xor data_in(174) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(179) xor data_in(180) xor data_in(187) xor data_in(192) xor data_in(193) xor data_in(194) xor data_in(197) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(204) xor data_in(210) xor data_in(211) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(223) xor data_in(224) xor data_in(225) xor data_in(227) xor data_in(229) xor data_in(231) xor data_in(233) xor data_in(234) xor data_in(237) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(242) xor data_in(244) xor data_in(247) xor data_in(248) xor data_in(251) xor data_in(252) xor data_in(254) xor data_in(255) xor data_in(256) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(264) xor data_in(265) xor data_in(267) xor data_in(270) xor data_in(273) xor data_in(274) xor data_in(275) xor data_in(277) xor data_in(278) xor data_in(279) xor data_in(281) xor data_in(282) xor data_in(283) xor data_in(285) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(296) xor data_in(297) xor data_in(303) xor data_in(304) xor data_in(308) xor data_in(309) xor data_in(310) xor data_in(313) xor data_in(314) xor data_in(315) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(324) xor data_in(325) xor data_in(330) xor data_in(331) xor data_in(334) xor data_in(335) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(340) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(350) xor data_in(351) xor data_in(354) xor data_in(356) xor data_in(358) xor data_in(360) xor data_in(361) xor data_in(364) xor data_in(366) xor data_in(368) xor data_in(370) xor data_in(371) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(379) xor data_in(382) xor data_in(387) xor data_in(389) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(398) xor data_in(400) xor data_in(401) xor data_in(402) xor data_in(403) xor data_in(404) xor data_in(406) xor data_in(407) xor data_in(408) xor data_in(411) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(418) xor data_in(421) xor data_in(423) xor data_in(424) xor data_in(426) xor data_in(427) xor data_in(430) xor data_in(431) xor data_in(434) xor data_in(436) xor data_in(438) xor data_in(439) xor data_in(442) xor data_in(447) xor data_in(448) xor data_in(451) xor data_in(452) xor data_in(454) xor data_in(457) xor data_in(461) xor data_in(462) xor data_in(464) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(470) xor data_in(471) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(482) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(500) xor data_in(501) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(509) xor data_in(510) xor data_in(511);
    crc_out(18) <= crc_in(0) xor crc_in(2) xor crc_in(3) xor crc_in(4) xor crc_in(5) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(10) xor crc_in(12) xor crc_in(16) xor crc_in(17) xor crc_in(18) xor crc_in(21) xor crc_in(22) xor crc_in(25) xor crc_in(26) xor crc_in(27) xor crc_in(29) xor crc_in(30) xor crc_in(35) xor crc_in(36) xor crc_in(40) xor crc_in(42) xor crc_in(43) xor crc_in(46) xor crc_in(47) xor crc_in(48) xor crc_in(51) xor crc_in(52) xor crc_in(55) xor crc_in(59) xor crc_in(61) xor data_in(0) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(12) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(21) xor data_in(22) xor data_in(25) xor data_in(26) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(35) xor data_in(36) xor data_in(40) xor data_in(42) xor data_in(43) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(52) xor data_in(55) xor data_in(59) xor data_in(61) xor data_in(64) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(75) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(85) xor data_in(86) xor data_in(88) xor data_in(89) xor data_in(90) xor data_in(95) xor data_in(96) xor data_in(102) xor data_in(106) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(112) xor data_in(115) xor data_in(117) xor data_in(118) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(125) xor data_in(126) xor data_in(130) xor data_in(132) xor data_in(138) xor data_in(139) xor data_in(141) xor data_in(142) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(154) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(158) xor data_in(160) xor data_in(162) xor data_in(163) xor data_in(166) xor data_in(179) xor data_in(180) xor data_in(182) xor data_in(184) xor data_in(186) xor data_in(188) xor data_in(190) xor data_in(193) xor data_in(195) xor data_in(197) xor data_in(198) xor data_in(201) xor data_in(202) xor data_in(204) xor data_in(206) xor data_in(207) xor data_in(208) xor data_in(214) xor data_in(216) xor data_in(218) xor data_in(221) xor data_in(222) xor data_in(229) xor data_in(231) xor data_in(233) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(243) xor data_in(248) xor data_in(249) xor data_in(253) xor data_in(254) xor data_in(255) xor data_in(256) xor data_in(257) xor data_in(258) xor data_in(260) xor data_in(261) xor data_in(263) xor data_in(264) xor data_in(265) xor data_in(267) xor data_in(269) xor data_in(271) xor data_in(274) xor data_in(279) xor data_in(280) xor data_in(281) xor data_in(282) xor data_in(283) xor data_in(284) xor data_in(286) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(292) xor data_in(295) xor data_in(299) xor data_in(300) xor data_in(302) xor data_in(303) xor data_in(305) xor data_in(310) xor data_in(311) xor data_in(313) xor data_in(315) xor data_in(316) xor data_in(319) xor data_in(322) xor data_in(324) xor data_in(327) xor data_in(330) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(341) xor data_in(343) xor data_in(344) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(351) xor data_in(353) xor data_in(356) xor data_in(358) xor data_in(359) xor data_in(361) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(368) xor data_in(369) xor data_in(371) xor data_in(373) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(382) xor data_in(383) xor data_in(385) xor data_in(387) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(396) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(402) xor data_in(403) xor data_in(404) xor data_in(407) xor data_in(413) xor data_in(415) xor data_in(420) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(425) xor data_in(427) xor data_in(428) xor data_in(429) xor data_in(430) xor data_in(432) xor data_in(434) xor data_in(437) xor data_in(438) xor data_in(440) xor data_in(442) xor data_in(443) xor data_in(448) xor data_in(454) xor data_in(455) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(472) xor data_in(474) xor data_in(476) xor data_in(479) xor data_in(480) xor data_in(483) xor data_in(484) xor data_in(486) xor data_in(489) xor data_in(491) xor data_in(494) xor data_in(495) xor data_in(498) xor data_in(499) xor data_in(501) xor data_in(502) xor data_in(503) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(509) xor data_in(511);
    crc_out(19) <= crc_in(1) xor crc_in(2) xor crc_in(3) xor crc_in(4) xor crc_in(6) xor crc_in(9) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(14) xor crc_in(15) xor crc_in(17) xor crc_in(18) xor crc_in(19) xor crc_in(21) xor crc_in(23) xor crc_in(24) xor crc_in(26) xor crc_in(27) xor crc_in(28) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(37) xor crc_in(44) xor crc_in(45) xor crc_in(48) xor crc_in(49) xor crc_in(50) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(6) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(37) xor data_in(44) xor data_in(45) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(65) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(73) xor data_in(77) xor data_in(78) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(85) xor data_in(89) xor data_in(90) xor data_in(91) xor data_in(92) xor data_in(95) xor data_in(96) xor data_in(97) xor data_in(102) xor data_in(104) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(114) xor data_in(116) xor data_in(118) xor data_in(120) xor data_in(121) xor data_in(127) xor data_in(129) xor data_in(130) xor data_in(131) xor data_in(132) xor data_in(133) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(141) xor data_in(144) xor data_in(145) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(154) xor data_in(159) xor data_in(160) xor data_in(161) xor data_in(163) xor data_in(165) xor data_in(166) xor data_in(168) xor data_in(170) xor data_in(171) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(182) xor data_in(183) xor data_in(184) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(189) xor data_in(190) xor data_in(191) xor data_in(196) xor data_in(197) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(202) xor data_in(203) xor data_in(204) xor data_in(206) xor data_in(209) xor data_in(211) xor data_in(212) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(222) xor data_in(224) xor data_in(225) xor data_in(226) xor data_in(228) xor data_in(229) xor data_in(231) xor data_in(233) xor data_in(235) xor data_in(236) xor data_in(238) xor data_in(240) xor data_in(241) xor data_in(244) xor data_in(245) xor data_in(249) xor data_in(250) xor data_in(252) xor data_in(255) xor data_in(256) xor data_in(257) xor data_in(259) xor data_in(261) xor data_in(263) xor data_in(265) xor data_in(267) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(276) xor data_in(278) xor data_in(280) xor data_in(282) xor data_in(283) xor data_in(284) xor data_in(285) xor data_in(289) xor data_in(290) xor data_in(293) xor data_in(295) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(301) xor data_in(302) xor data_in(306) xor data_in(309) xor data_in(311) xor data_in(312) xor data_in(313) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(326) xor data_in(327) xor data_in(328) xor data_in(330) xor data_in(332) xor data_in(333) xor data_in(335) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(342) xor data_in(343) xor data_in(346) xor data_in(350) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(363) xor data_in(365) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(373) xor data_in(374) xor data_in(377) xor data_in(378) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(385) xor data_in(386) xor data_in(387) xor data_in(394) xor data_in(395) xor data_in(398) xor data_in(399) xor data_in(401) xor data_in(402) xor data_in(403) xor data_in(404) xor data_in(409) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(417) xor data_in(419) xor data_in(420) xor data_in(422) xor data_in(426) xor data_in(428) xor data_in(433) xor data_in(434) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(456) xor data_in(463) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(473) xor data_in(474) xor data_in(478) xor data_in(480) xor data_in(481) xor data_in(485) xor data_in(486) xor data_in(488) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(495) xor data_in(498) xor data_in(500) xor data_in(502) xor data_in(506) xor data_in(507);
    crc_out(20) <= crc_in(0) xor crc_in(2) xor crc_in(3) xor crc_in(4) xor crc_in(5) xor crc_in(7) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(15) xor crc_in(16) xor crc_in(18) xor crc_in(19) xor crc_in(20) xor crc_in(22) xor crc_in(24) xor crc_in(25) xor crc_in(27) xor crc_in(28) xor crc_in(29) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(38) xor crc_in(45) xor crc_in(46) xor crc_in(49) xor crc_in(50) xor crc_in(51) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor data_in(0) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(38) xor data_in(45) xor data_in(46) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(66) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(74) xor data_in(78) xor data_in(79) xor data_in(82) xor data_in(83) xor data_in(84) xor data_in(86) xor data_in(90) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(96) xor data_in(97) xor data_in(98) xor data_in(103) xor data_in(105) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(115) xor data_in(117) xor data_in(119) xor data_in(121) xor data_in(122) xor data_in(128) xor data_in(130) xor data_in(131) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(142) xor data_in(145) xor data_in(146) xor data_in(149) xor data_in(150) xor data_in(152) xor data_in(155) xor data_in(160) xor data_in(161) xor data_in(162) xor data_in(164) xor data_in(166) xor data_in(167) xor data_in(169) xor data_in(171) xor data_in(172) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(183) xor data_in(184) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(190) xor data_in(191) xor data_in(192) xor data_in(197) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(203) xor data_in(204) xor data_in(205) xor data_in(207) xor data_in(210) xor data_in(212) xor data_in(213) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(223) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(229) xor data_in(230) xor data_in(232) xor data_in(234) xor data_in(236) xor data_in(237) xor data_in(239) xor data_in(241) xor data_in(242) xor data_in(245) xor data_in(246) xor data_in(250) xor data_in(251) xor data_in(253) xor data_in(256) xor data_in(257) xor data_in(258) xor data_in(260) xor data_in(262) xor data_in(264) xor data_in(266) xor data_in(268) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(277) xor data_in(279) xor data_in(281) xor data_in(283) xor data_in(284) xor data_in(285) xor data_in(286) xor data_in(290) xor data_in(291) xor data_in(294) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(302) xor data_in(303) xor data_in(307) xor data_in(310) xor data_in(312) xor data_in(313) xor data_in(314) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(327) xor data_in(328) xor data_in(329) xor data_in(331) xor data_in(333) xor data_in(334) xor data_in(336) xor data_in(337) xor data_in(338) xor data_in(340) xor data_in(343) xor data_in(344) xor data_in(347) xor data_in(351) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(364) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(374) xor data_in(375) xor data_in(378) xor data_in(379) xor data_in(383) xor data_in(384) xor data_in(385) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(395) xor data_in(396) xor data_in(399) xor data_in(400) xor data_in(402) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(410) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(418) xor data_in(420) xor data_in(421) xor data_in(423) xor data_in(427) xor data_in(429) xor data_in(434) xor data_in(435) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(456) xor data_in(457) xor data_in(464) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(474) xor data_in(475) xor data_in(479) xor data_in(481) xor data_in(482) xor data_in(486) xor data_in(487) xor data_in(489) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(496) xor data_in(499) xor data_in(501) xor data_in(503) xor data_in(507) xor data_in(508);
    crc_out(21) <= crc_in(1) xor crc_in(3) xor crc_in(4) xor crc_in(5) xor crc_in(6) xor crc_in(8) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(16) xor crc_in(17) xor crc_in(19) xor crc_in(20) xor crc_in(21) xor crc_in(23) xor crc_in(25) xor crc_in(26) xor crc_in(28) xor crc_in(29) xor crc_in(30) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(39) xor crc_in(46) xor crc_in(47) xor crc_in(50) xor crc_in(51) xor crc_in(52) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(8) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(39) xor data_in(46) xor data_in(47) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(67) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(75) xor data_in(79) xor data_in(80) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(87) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(94) xor data_in(97) xor data_in(98) xor data_in(99) xor data_in(104) xor data_in(106) xor data_in(109) xor data_in(110) xor data_in(111) xor data_in(116) xor data_in(118) xor data_in(120) xor data_in(122) xor data_in(123) xor data_in(129) xor data_in(131) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(138) xor data_in(139) xor data_in(140) xor data_in(143) xor data_in(146) xor data_in(147) xor data_in(150) xor data_in(151) xor data_in(153) xor data_in(156) xor data_in(161) xor data_in(162) xor data_in(163) xor data_in(165) xor data_in(167) xor data_in(168) xor data_in(170) xor data_in(172) xor data_in(173) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(184) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(191) xor data_in(192) xor data_in(193) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(204) xor data_in(205) xor data_in(206) xor data_in(208) xor data_in(211) xor data_in(213) xor data_in(214) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(224) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(230) xor data_in(231) xor data_in(233) xor data_in(235) xor data_in(237) xor data_in(238) xor data_in(240) xor data_in(242) xor data_in(243) xor data_in(246) xor data_in(247) xor data_in(251) xor data_in(252) xor data_in(254) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(261) xor data_in(263) xor data_in(265) xor data_in(267) xor data_in(269) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(278) xor data_in(280) xor data_in(282) xor data_in(284) xor data_in(285) xor data_in(286) xor data_in(287) xor data_in(291) xor data_in(292) xor data_in(295) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(303) xor data_in(304) xor data_in(308) xor data_in(311) xor data_in(313) xor data_in(314) xor data_in(315) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(328) xor data_in(329) xor data_in(330) xor data_in(332) xor data_in(334) xor data_in(335) xor data_in(337) xor data_in(338) xor data_in(339) xor data_in(341) xor data_in(344) xor data_in(345) xor data_in(348) xor data_in(352) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(360) xor data_in(361) xor data_in(362) xor data_in(365) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(375) xor data_in(376) xor data_in(379) xor data_in(380) xor data_in(384) xor data_in(385) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(396) xor data_in(397) xor data_in(400) xor data_in(401) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(411) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(419) xor data_in(421) xor data_in(422) xor data_in(424) xor data_in(428) xor data_in(430) xor data_in(435) xor data_in(436) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(454) xor data_in(455) xor data_in(456) xor data_in(457) xor data_in(458) xor data_in(465) xor data_in(469) xor data_in(470) xor data_in(471) xor data_in(475) xor data_in(476) xor data_in(480) xor data_in(482) xor data_in(483) xor data_in(487) xor data_in(488) xor data_in(490) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(497) xor data_in(500) xor data_in(502) xor data_in(504) xor data_in(508) xor data_in(509);
    crc_out(22) <= crc_in(0) xor crc_in(2) xor crc_in(4) xor crc_in(5) xor crc_in(6) xor crc_in(7) xor crc_in(9) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(17) xor crc_in(18) xor crc_in(20) xor crc_in(21) xor crc_in(22) xor crc_in(24) xor crc_in(26) xor crc_in(27) xor crc_in(29) xor crc_in(30) xor crc_in(31) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(40) xor crc_in(47) xor crc_in(48) xor crc_in(51) xor crc_in(52) xor crc_in(53) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(40) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(68) xor data_in(72) xor data_in(73) xor data_in(74) xor data_in(76) xor data_in(80) xor data_in(81) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(88) xor data_in(92) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(98) xor data_in(99) xor data_in(100) xor data_in(105) xor data_in(107) xor data_in(110) xor data_in(111) xor data_in(112) xor data_in(117) xor data_in(119) xor data_in(121) xor data_in(123) xor data_in(124) xor data_in(130) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(136) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(144) xor data_in(147) xor data_in(148) xor data_in(151) xor data_in(152) xor data_in(154) xor data_in(157) xor data_in(162) xor data_in(163) xor data_in(164) xor data_in(166) xor data_in(168) xor data_in(169) xor data_in(171) xor data_in(173) xor data_in(174) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(183) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(190) xor data_in(192) xor data_in(193) xor data_in(194) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(209) xor data_in(212) xor data_in(214) xor data_in(215) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(225) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(231) xor data_in(232) xor data_in(234) xor data_in(236) xor data_in(238) xor data_in(239) xor data_in(241) xor data_in(243) xor data_in(244) xor data_in(247) xor data_in(248) xor data_in(252) xor data_in(253) xor data_in(255) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(262) xor data_in(264) xor data_in(266) xor data_in(268) xor data_in(270) xor data_in(272) xor data_in(273) xor data_in(275) xor data_in(279) xor data_in(281) xor data_in(283) xor data_in(285) xor data_in(286) xor data_in(287) xor data_in(288) xor data_in(292) xor data_in(293) xor data_in(296) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(304) xor data_in(305) xor data_in(309) xor data_in(312) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(319) xor data_in(320) xor data_in(321) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(333) xor data_in(335) xor data_in(336) xor data_in(338) xor data_in(339) xor data_in(340) xor data_in(342) xor data_in(345) xor data_in(346) xor data_in(349) xor data_in(353) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(361) xor data_in(362) xor data_in(363) xor data_in(366) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(376) xor data_in(377) xor data_in(380) xor data_in(381) xor data_in(385) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(397) xor data_in(398) xor data_in(401) xor data_in(402) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(407) xor data_in(412) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(420) xor data_in(422) xor data_in(423) xor data_in(425) xor data_in(429) xor data_in(431) xor data_in(436) xor data_in(437) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(455) xor data_in(456) xor data_in(457) xor data_in(458) xor data_in(459) xor data_in(466) xor data_in(470) xor data_in(471) xor data_in(472) xor data_in(476) xor data_in(477) xor data_in(481) xor data_in(483) xor data_in(484) xor data_in(488) xor data_in(489) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(498) xor data_in(501) xor data_in(503) xor data_in(505) xor data_in(509) xor data_in(510);
    crc_out(23) <= crc_in(0) xor crc_in(1) xor crc_in(3) xor crc_in(5) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(10) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(18) xor crc_in(19) xor crc_in(21) xor crc_in(22) xor crc_in(23) xor crc_in(25) xor crc_in(27) xor crc_in(28) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(41) xor crc_in(48) xor crc_in(49) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(41) xor data_in(48) xor data_in(49) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(62) xor data_in(63) xor data_in(64) xor data_in(69) xor data_in(73) xor data_in(74) xor data_in(75) xor data_in(77) xor data_in(81) xor data_in(82) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(89) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(99) xor data_in(100) xor data_in(101) xor data_in(106) xor data_in(108) xor data_in(111) xor data_in(112) xor data_in(113) xor data_in(118) xor data_in(120) xor data_in(122) xor data_in(124) xor data_in(125) xor data_in(131) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(140) xor data_in(141) xor data_in(142) xor data_in(145) xor data_in(148) xor data_in(149) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(158) xor data_in(163) xor data_in(164) xor data_in(165) xor data_in(167) xor data_in(169) xor data_in(170) xor data_in(172) xor data_in(174) xor data_in(175) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(183) xor data_in(184) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(190) xor data_in(191) xor data_in(193) xor data_in(194) xor data_in(195) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(204) xor data_in(206) xor data_in(207) xor data_in(208) xor data_in(210) xor data_in(213) xor data_in(215) xor data_in(216) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(223) xor data_in(226) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(232) xor data_in(233) xor data_in(235) xor data_in(237) xor data_in(239) xor data_in(240) xor data_in(242) xor data_in(244) xor data_in(245) xor data_in(248) xor data_in(249) xor data_in(253) xor data_in(254) xor data_in(256) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(263) xor data_in(265) xor data_in(267) xor data_in(269) xor data_in(271) xor data_in(273) xor data_in(274) xor data_in(276) xor data_in(280) xor data_in(282) xor data_in(284) xor data_in(286) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(293) xor data_in(294) xor data_in(297) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(305) xor data_in(306) xor data_in(310) xor data_in(313) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(334) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(340) xor data_in(341) xor data_in(343) xor data_in(346) xor data_in(347) xor data_in(350) xor data_in(354) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(362) xor data_in(363) xor data_in(364) xor data_in(367) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(377) xor data_in(378) xor data_in(381) xor data_in(382) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(398) xor data_in(399) xor data_in(402) xor data_in(403) xor data_in(405) xor data_in(406) xor data_in(407) xor data_in(408) xor data_in(413) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(421) xor data_in(423) xor data_in(424) xor data_in(426) xor data_in(430) xor data_in(432) xor data_in(437) xor data_in(438) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(456) xor data_in(457) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(467) xor data_in(471) xor data_in(472) xor data_in(473) xor data_in(477) xor data_in(478) xor data_in(482) xor data_in(484) xor data_in(485) xor data_in(489) xor data_in(490) xor data_in(492) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(497) xor data_in(499) xor data_in(502) xor data_in(504) xor data_in(506) xor data_in(510) xor data_in(511);
    crc_out(24) <= crc_in(0) xor crc_in(1) xor crc_in(4) xor crc_in(5) xor crc_in(6) xor crc_in(9) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(16) xor crc_in(17) xor crc_in(19) xor crc_in(20) xor crc_in(21) xor crc_in(23) xor crc_in(26) xor crc_in(28) xor crc_in(29) xor crc_in(31) xor crc_in(33) xor crc_in(35) xor crc_in(37) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(45) xor crc_in(47) xor crc_in(49) xor crc_in(52) xor crc_in(58) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(33) xor data_in(35) xor data_in(37) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(45) xor data_in(47) xor data_in(49) xor data_in(52) xor data_in(58) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(64) xor data_in(65) xor data_in(69) xor data_in(71) xor data_in(72) xor data_in(75) xor data_in(77) xor data_in(79) xor data_in(80) xor data_in(85) xor data_in(88) xor data_in(90) xor data_in(92) xor data_in(94) xor data_in(96) xor data_in(97) xor data_in(100) xor data_in(101) xor data_in(103) xor data_in(104) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(111) xor data_in(112) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(124) xor data_in(125) xor data_in(129) xor data_in(130) xor data_in(134) xor data_in(135) xor data_in(139) xor data_in(140) xor data_in(149) xor data_in(151) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(157) xor data_in(158) xor data_in(159) xor data_in(160) xor data_in(167) xor data_in(173) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(183) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(191) xor data_in(192) xor data_in(195) xor data_in(196) xor data_in(197) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(206) xor data_in(209) xor data_in(212) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(232) xor data_in(235) xor data_in(237) xor data_in(238) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(242) xor data_in(243) xor data_in(246) xor data_in(249) xor data_in(250) xor data_in(252) xor data_in(255) xor data_in(257) xor data_in(258) xor data_in(260) xor data_in(261) xor data_in(263) xor data_in(267) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(274) xor data_in(276) xor data_in(277) xor data_in(278) xor data_in(283) xor data_in(285) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(294) xor data_in(297) xor data_in(299) xor data_in(301) xor data_in(306) xor data_in(307) xor data_in(309) xor data_in(311) xor data_in(313) xor data_in(316) xor data_in(317) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(330) xor data_in(334) xor data_in(335) xor data_in(337) xor data_in(339) xor data_in(341) xor data_in(342) xor data_in(343) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(349) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(356) xor data_in(357) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(362) xor data_in(365) xor data_in(367) xor data_in(370) xor data_in(371) xor data_in(374) xor data_in(375) xor data_in(378) xor data_in(380) xor data_in(383) xor data_in(385) xor data_in(389) xor data_in(390) xor data_in(393) xor data_in(395) xor data_in(397) xor data_in(398) xor data_in(399) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(407) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(416) xor data_in(418) xor data_in(420) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(425) xor data_in(427) xor data_in(429) xor data_in(430) xor data_in(433) xor data_in(434) xor data_in(435) xor data_in(442) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(457) xor data_in(458) xor data_in(462) xor data_in(463) xor data_in(466) xor data_in(468) xor data_in(470) xor data_in(471) xor data_in(472) xor data_in(473) xor data_in(475) xor data_in(477) xor data_in(479) xor data_in(483) xor data_in(484) xor data_in(485) xor data_in(487) xor data_in(488) xor data_in(490) xor data_in(495) xor data_in(497) xor data_in(499) xor data_in(500) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(510) xor data_in(511);
    crc_out(25) <= crc_in(1) xor crc_in(6) xor crc_in(8) xor crc_in(11) xor crc_in(15) xor crc_in(17) xor crc_in(18) xor crc_in(20) xor crc_in(27) xor crc_in(29) xor crc_in(30) xor crc_in(34) xor crc_in(38) xor crc_in(41) xor crc_in(42) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(47) xor crc_in(48) xor crc_in(52) xor crc_in(54) xor crc_in(55) xor crc_in(58) xor crc_in(61) xor crc_in(63) xor data_in(1) xor data_in(6) xor data_in(8) xor data_in(11) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(34) xor data_in(38) xor data_in(41) xor data_in(42) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(52) xor data_in(54) xor data_in(55) xor data_in(58) xor data_in(61) xor data_in(63) xor data_in(64) xor data_in(65) xor data_in(66) xor data_in(69) xor data_in(71) xor data_in(73) xor data_in(74) xor data_in(77) xor data_in(79) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(85) xor data_in(87) xor data_in(89) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(97) xor data_in(98) xor data_in(101) xor data_in(103) xor data_in(105) xor data_in(109) xor data_in(112) xor data_in(114) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(124) xor data_in(125) xor data_in(129) xor data_in(131) xor data_in(132) xor data_in(135) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(142) xor data_in(143) xor data_in(146) xor data_in(151) xor data_in(153) xor data_in(155) xor data_in(157) xor data_in(159) xor data_in(161) xor data_in(164) xor data_in(165) xor data_in(166) xor data_in(167) xor data_in(170) xor data_in(171) xor data_in(174) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(180) xor data_in(182) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(192) xor data_in(193) xor data_in(194) xor data_in(196) xor data_in(198) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(206) xor data_in(208) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(216) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(224) xor data_in(225) xor data_in(227) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(234) xor data_in(235) xor data_in(237) xor data_in(238) xor data_in(240) xor data_in(241) xor data_in(243) xor data_in(244) xor data_in(245) xor data_in(247) xor data_in(250) xor data_in(251) xor data_in(252) xor data_in(253) xor data_in(254) xor data_in(256) xor data_in(259) xor data_in(261) xor data_in(263) xor data_in(266) xor data_in(267) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(276) xor data_in(277) xor data_in(279) xor data_in(281) xor data_in(284) xor data_in(286) xor data_in(287) xor data_in(288) xor data_in(290) xor data_in(292) xor data_in(297) xor data_in(299) xor data_in(303) xor data_in(304) xor data_in(307) xor data_in(308) xor data_in(309) xor data_in(310) xor data_in(312) xor data_in(313) xor data_in(317) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(325) xor data_in(328) xor data_in(330) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(336) xor data_in(339) xor data_in(342) xor data_in(345) xor data_in(347) xor data_in(349) xor data_in(350) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(360) xor data_in(361) xor data_in(364) xor data_in(366) xor data_in(367) xor data_in(371) xor data_in(373) xor data_in(375) xor data_in(376) xor data_in(380) xor data_in(381) xor data_in(382) xor data_in(384) xor data_in(385) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(390) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(399) xor data_in(404) xor data_in(406) xor data_in(407) xor data_in(409) xor data_in(412) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(420) xor data_in(422) xor data_in(426) xor data_in(428) xor data_in(429) xor data_in(436) xor data_in(438) xor data_in(439) xor data_in(442) xor data_in(443) xor data_in(447) xor data_in(448) xor data_in(452) xor data_in(455) xor data_in(458) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(464) xor data_in(466) xor data_in(467) xor data_in(469) xor data_in(470) xor data_in(472) xor data_in(473) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(480) xor data_in(485) xor data_in(487) xor data_in(489) xor data_in(493) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(503) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(509) xor data_in(510) xor data_in(511);
    crc_out(26) <= crc_in(0) xor crc_in(5) xor crc_in(8) xor crc_in(9) xor crc_in(10) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(18) xor crc_in(19) xor crc_in(22) xor crc_in(24) xor crc_in(28) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(35) xor crc_in(36) xor crc_in(39) xor crc_in(41) xor crc_in(42) xor crc_in(46) xor crc_in(48) xor crc_in(49) xor crc_in(50) xor crc_in(52) xor crc_in(54) xor crc_in(56) xor crc_in(58) xor data_in(0) xor data_in(5) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(22) xor data_in(24) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(35) xor data_in(36) xor data_in(39) xor data_in(41) xor data_in(42) xor data_in(46) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(52) xor data_in(54) xor data_in(56) xor data_in(58) xor data_in(64) xor data_in(65) xor data_in(66) xor data_in(67) xor data_in(69) xor data_in(71) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(79) xor data_in(84) xor data_in(85) xor data_in(87) xor data_in(88) xor data_in(90) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(98) xor data_in(99) xor data_in(103) xor data_in(106) xor data_in(108) xor data_in(111) xor data_in(114) xor data_in(115) xor data_in(119) xor data_in(121) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(129) xor data_in(133) xor data_in(137) xor data_in(141) xor data_in(142) xor data_in(144) xor data_in(146) xor data_in(147) xor data_in(150) xor data_in(151) xor data_in(155) xor data_in(157) xor data_in(162) xor data_in(164) xor data_in(170) xor data_in(172) xor data_in(179) xor data_in(182) xor data_in(183) xor data_in(184) xor data_in(186) xor data_in(188) xor data_in(189) xor data_in(193) xor data_in(195) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(208) xor data_in(209) xor data_in(213) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(224) xor data_in(229) xor data_in(230) xor data_in(234) xor data_in(237) xor data_in(238) xor data_in(241) xor data_in(244) xor data_in(246) xor data_in(248) xor data_in(251) xor data_in(253) xor data_in(255) xor data_in(257) xor data_in(258) xor data_in(260) xor data_in(263) xor data_in(266) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(275) xor data_in(276) xor data_in(277) xor data_in(280) xor data_in(281) xor data_in(282) xor data_in(285) xor data_in(289) xor data_in(293) xor data_in(295) xor data_in(297) xor data_in(299) xor data_in(302) xor data_in(303) xor data_in(305) xor data_in(308) xor data_in(310) xor data_in(311) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(325) xor data_in(327) xor data_in(329) xor data_in(330) xor data_in(332) xor data_in(335) xor data_in(336) xor data_in(337) xor data_in(338) xor data_in(339) xor data_in(344) xor data_in(345) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(358) xor data_in(361) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(373) xor data_in(374) xor data_in(376) xor data_in(377) xor data_in(379) xor data_in(380) xor data_in(381) xor data_in(383) xor data_in(386) xor data_in(389) xor data_in(392) xor data_in(394) xor data_in(396) xor data_in(407) xor data_in(409) xor data_in(410) xor data_in(412) xor data_in(415) xor data_in(419) xor data_in(420) xor data_in(424) xor data_in(427) xor data_in(431) xor data_in(434) xor data_in(435) xor data_in(437) xor data_in(438) xor data_in(440) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(448) xor data_in(452) xor data_in(454) xor data_in(456) xor data_in(460) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(473) xor data_in(475) xor data_in(476) xor data_in(481) xor data_in(484) xor data_in(487) xor data_in(490) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(496) xor data_in(498) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(503) xor data_in(506) xor data_in(507) xor data_in(511);
    crc_out(27) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(5) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(16) xor crc_in(17) xor crc_in(19) xor crc_in(20) xor crc_in(21) xor crc_in(22) xor crc_in(23) xor crc_in(24) xor crc_in(25) xor crc_in(29) xor crc_in(31) xor crc_in(33) xor crc_in(37) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(45) xor crc_in(49) xor crc_in(51) xor crc_in(52) xor crc_in(54) xor crc_in(57) xor crc_in(58) xor crc_in(62) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(29) xor data_in(31) xor data_in(33) xor data_in(37) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(45) xor data_in(49) xor data_in(51) xor data_in(52) xor data_in(54) xor data_in(57) xor data_in(58) xor data_in(62) xor data_in(65) xor data_in(66) xor data_in(67) xor data_in(68) xor data_in(69) xor data_in(71) xor data_in(74) xor data_in(79) xor data_in(82) xor data_in(83) xor data_in(87) xor data_in(88) xor data_in(89) xor data_in(91) xor data_in(92) xor data_in(94) xor data_in(96) xor data_in(99) xor data_in(100) xor data_in(102) xor data_in(103) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(111) xor data_in(112) xor data_in(113) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(119) xor data_in(123) xor data_in(125) xor data_in(129) xor data_in(132) xor data_in(134) xor data_in(136) xor data_in(137) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(145) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(150) xor data_in(154) xor data_in(155) xor data_in(157) xor data_in(160) xor data_in(163) xor data_in(164) xor data_in(166) xor data_in(167) xor data_in(168) xor data_in(170) xor data_in(173) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(183) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(189) xor data_in(196) xor data_in(197) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(207) xor data_in(208) xor data_in(209) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(217) xor data_in(219) xor data_in(221) xor data_in(222) xor data_in(224) xor data_in(226) xor data_in(228) xor data_in(229) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(247) xor data_in(249) xor data_in(256) xor data_in(259) xor data_in(261) xor data_in(262) xor data_in(263) xor data_in(266) xor data_in(268) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(277) xor data_in(282) xor data_in(283) xor data_in(286) xor data_in(287) xor data_in(288) xor data_in(290) xor data_in(291) xor data_in(294) xor data_in(295) xor data_in(296) xor data_in(297) xor data_in(299) xor data_in(302) xor data_in(306) xor data_in(311) xor data_in(312) xor data_in(313) xor data_in(314) xor data_in(318) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(325) xor data_in(327) xor data_in(328) xor data_in(332) xor data_in(334) xor data_in(336) xor data_in(337) xor data_in(343) xor data_in(344) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(363) xor data_in(365) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(381) xor data_in(384) xor data_in(385) xor data_in(388) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(398) xor data_in(400) xor data_in(405) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(417) xor data_in(419) xor data_in(423) xor data_in(424) xor data_in(425) xor data_in(428) xor data_in(429) xor data_in(430) xor data_in(431) xor data_in(432) xor data_in(434) xor data_in(436) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(452) xor data_in(454) xor data_in(455) xor data_in(457) xor data_in(459) xor data_in(460) xor data_in(462) xor data_in(463) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(471) xor data_in(475) xor data_in(476) xor data_in(478) xor data_in(482) xor data_in(484) xor data_in(485) xor data_in(486) xor data_in(487) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(497) xor data_in(498) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(510);
    crc_out(28) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(3) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(10) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(17) xor crc_in(18) xor crc_in(20) xor crc_in(21) xor crc_in(22) xor crc_in(23) xor crc_in(24) xor crc_in(25) xor crc_in(26) xor crc_in(30) xor crc_in(32) xor crc_in(34) xor crc_in(38) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(46) xor crc_in(50) xor crc_in(52) xor crc_in(53) xor crc_in(55) xor crc_in(58) xor crc_in(59) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(30) xor data_in(32) xor data_in(34) xor data_in(38) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(46) xor data_in(50) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(58) xor data_in(59) xor data_in(63) xor data_in(66) xor data_in(67) xor data_in(68) xor data_in(69) xor data_in(70) xor data_in(72) xor data_in(75) xor data_in(80) xor data_in(83) xor data_in(84) xor data_in(88) xor data_in(89) xor data_in(90) xor data_in(92) xor data_in(93) xor data_in(95) xor data_in(97) xor data_in(100) xor data_in(101) xor data_in(103) xor data_in(104) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(111) xor data_in(112) xor data_in(113) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(120) xor data_in(124) xor data_in(126) xor data_in(130) xor data_in(133) xor data_in(135) xor data_in(137) xor data_in(138) xor data_in(140) xor data_in(141) xor data_in(142) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(155) xor data_in(156) xor data_in(158) xor data_in(161) xor data_in(164) xor data_in(165) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(171) xor data_in(174) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(183) xor data_in(184) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(190) xor data_in(197) xor data_in(198) xor data_in(202) xor data_in(203) xor data_in(204) xor data_in(206) xor data_in(208) xor data_in(209) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(218) xor data_in(220) xor data_in(222) xor data_in(223) xor data_in(225) xor data_in(227) xor data_in(229) xor data_in(230) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(237) xor data_in(238) xor data_in(239) xor data_in(248) xor data_in(250) xor data_in(257) xor data_in(260) xor data_in(262) xor data_in(263) xor data_in(264) xor data_in(267) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(278) xor data_in(283) xor data_in(284) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(291) xor data_in(292) xor data_in(295) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(300) xor data_in(303) xor data_in(307) xor data_in(312) xor data_in(313) xor data_in(314) xor data_in(315) xor data_in(319) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(326) xor data_in(328) xor data_in(329) xor data_in(333) xor data_in(335) xor data_in(337) xor data_in(338) xor data_in(344) xor data_in(345) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(364) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(378) xor data_in(379) xor data_in(380) xor data_in(382) xor data_in(385) xor data_in(386) xor data_in(389) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(399) xor data_in(401) xor data_in(406) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(418) xor data_in(420) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(429) xor data_in(430) xor data_in(431) xor data_in(432) xor data_in(433) xor data_in(435) xor data_in(437) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(453) xor data_in(455) xor data_in(456) xor data_in(458) xor data_in(460) xor data_in(461) xor data_in(463) xor data_in(464) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(471) xor data_in(472) xor data_in(476) xor data_in(477) xor data_in(479) xor data_in(483) xor data_in(485) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(497) xor data_in(498) xor data_in(499) xor data_in(501) xor data_in(502) xor data_in(503) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(511);
    crc_out(29) <= crc_in(1) xor crc_in(3) xor crc_in(4) xor crc_in(5) xor crc_in(9) xor crc_in(11) xor crc_in(12) xor crc_in(18) xor crc_in(19) xor crc_in(23) xor crc_in(25) xor crc_in(26) xor crc_in(27) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(35) xor crc_in(36) xor crc_in(39) xor crc_in(41) xor crc_in(42) xor crc_in(44) xor crc_in(45) xor crc_in(50) xor crc_in(51) xor crc_in(52) xor crc_in(55) xor crc_in(56) xor crc_in(58) xor crc_in(60) xor crc_in(62) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(18) xor data_in(19) xor data_in(23) xor data_in(25) xor data_in(26) xor data_in(27) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(35) xor data_in(36) xor data_in(39) xor data_in(41) xor data_in(42) xor data_in(44) xor data_in(45) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(55) xor data_in(56) xor data_in(58) xor data_in(60) xor data_in(62) xor data_in(64) xor data_in(67) xor data_in(68) xor data_in(72) xor data_in(73) xor data_in(74) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(84) xor data_in(86) xor data_in(87) xor data_in(89) xor data_in(90) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(98) xor data_in(101) xor data_in(103) xor data_in(105) xor data_in(108) xor data_in(109) xor data_in(112) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(129) xor data_in(130) xor data_in(131) xor data_in(132) xor data_in(134) xor data_in(137) xor data_in(140) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(154) xor data_in(155) xor data_in(158) xor data_in(159) xor data_in(160) xor data_in(162) xor data_in(164) xor data_in(167) xor data_in(169) xor data_in(171) xor data_in(172) xor data_in(176) xor data_in(180) xor data_in(183) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(190) xor data_in(191) xor data_in(194) xor data_in(197) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(203) xor data_in(206) xor data_in(208) xor data_in(209) xor data_in(210) xor data_in(213) xor data_in(216) xor data_in(218) xor data_in(219) xor data_in(221) xor data_in(225) xor data_in(229) xor data_in(232) xor data_in(233) xor data_in(237) xor data_in(238) xor data_in(240) xor data_in(242) xor data_in(245) xor data_in(249) xor data_in(251) xor data_in(252) xor data_in(254) xor data_in(261) xor data_in(262) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(276) xor data_in(278) xor data_in(279) xor data_in(281) xor data_in(284) xor data_in(285) xor data_in(287) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(295) xor data_in(296) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(308) xor data_in(309) xor data_in(315) xor data_in(316) xor data_in(318) xor data_in(322) xor data_in(324) xor data_in(325) xor data_in(326) xor data_in(329) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(336) xor data_in(340) xor data_in(343) xor data_in(344) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(355) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(362) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(369) xor data_in(370) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(385) xor data_in(386) xor data_in(388) xor data_in(390) xor data_in(391) xor data_in(394) xor data_in(395) xor data_in(397) xor data_in(398) xor data_in(402) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(411) xor data_in(414) xor data_in(416) xor data_in(417) xor data_in(420) xor data_in(423) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(429) xor data_in(432) xor data_in(433) xor data_in(435) xor data_in(436) xor data_in(439) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(449) xor data_in(452) xor data_in(453) xor data_in(456) xor data_in(457) xor data_in(460) xor data_in(463) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(469) xor data_in(472) xor data_in(473) xor data_in(474) xor data_in(475) xor data_in(480) xor data_in(489) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(497) xor data_in(500) xor data_in(502) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(509) xor data_in(510);
    crc_out(30) <= crc_in(2) xor crc_in(4) xor crc_in(5) xor crc_in(6) xor crc_in(10) xor crc_in(12) xor crc_in(13) xor crc_in(19) xor crc_in(20) xor crc_in(24) xor crc_in(26) xor crc_in(27) xor crc_in(28) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(36) xor crc_in(37) xor crc_in(40) xor crc_in(42) xor crc_in(43) xor crc_in(45) xor crc_in(46) xor crc_in(51) xor crc_in(52) xor crc_in(53) xor crc_in(56) xor crc_in(57) xor crc_in(59) xor crc_in(61) xor crc_in(63) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(19) xor data_in(20) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(36) xor data_in(37) xor data_in(40) xor data_in(42) xor data_in(43) xor data_in(45) xor data_in(46) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(56) xor data_in(57) xor data_in(59) xor data_in(61) xor data_in(63) xor data_in(65) xor data_in(68) xor data_in(69) xor data_in(73) xor data_in(74) xor data_in(75) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(87) xor data_in(88) xor data_in(90) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(97) xor data_in(99) xor data_in(102) xor data_in(104) xor data_in(106) xor data_in(109) xor data_in(110) xor data_in(113) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(128) xor data_in(130) xor data_in(131) xor data_in(132) xor data_in(133) xor data_in(135) xor data_in(138) xor data_in(141) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(150) xor data_in(152) xor data_in(155) xor data_in(156) xor data_in(159) xor data_in(160) xor data_in(161) xor data_in(163) xor data_in(165) xor data_in(168) xor data_in(170) xor data_in(172) xor data_in(173) xor data_in(177) xor data_in(181) xor data_in(184) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(190) xor data_in(191) xor data_in(192) xor data_in(195) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(204) xor data_in(207) xor data_in(209) xor data_in(210) xor data_in(211) xor data_in(214) xor data_in(217) xor data_in(219) xor data_in(220) xor data_in(222) xor data_in(226) xor data_in(230) xor data_in(233) xor data_in(234) xor data_in(238) xor data_in(239) xor data_in(241) xor data_in(243) xor data_in(246) xor data_in(250) xor data_in(252) xor data_in(253) xor data_in(255) xor data_in(262) xor data_in(263) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(275) xor data_in(277) xor data_in(279) xor data_in(280) xor data_in(282) xor data_in(285) xor data_in(286) xor data_in(288) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(296) xor data_in(297) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(304) xor data_in(309) xor data_in(310) xor data_in(316) xor data_in(317) xor data_in(319) xor data_in(323) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(330) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(337) xor data_in(341) xor data_in(344) xor data_in(345) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(356) xor data_in(360) xor data_in(361) xor data_in(362) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(366) xor data_in(370) xor data_in(371) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(386) xor data_in(387) xor data_in(389) xor data_in(391) xor data_in(392) xor data_in(395) xor data_in(396) xor data_in(398) xor data_in(399) xor data_in(403) xor data_in(406) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(412) xor data_in(415) xor data_in(417) xor data_in(418) xor data_in(421) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(430) xor data_in(433) xor data_in(434) xor data_in(436) xor data_in(437) xor data_in(440) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(450) xor data_in(453) xor data_in(454) xor data_in(457) xor data_in(458) xor data_in(461) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(470) xor data_in(473) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(481) xor data_in(490) xor data_in(492) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(498) xor data_in(501) xor data_in(503) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(510) xor data_in(511);
    crc_out(31) <= crc_in(0) xor crc_in(2) xor crc_in(3) xor crc_in(6) xor crc_in(8) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(15) xor crc_in(20) xor crc_in(22) xor crc_in(24) xor crc_in(25) xor crc_in(27) xor crc_in(28) xor crc_in(29) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(37) xor crc_in(38) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(50) xor crc_in(55) xor crc_in(57) xor crc_in(59) xor crc_in(60) xor data_in(0) xor data_in(2) xor data_in(3) xor data_in(6) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(15) xor data_in(20) xor data_in(22) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(50) xor data_in(55) xor data_in(57) xor data_in(59) xor data_in(60) xor data_in(64) xor data_in(66) xor data_in(71) xor data_in(72) xor data_in(75) xor data_in(77) xor data_in(78) xor data_in(81) xor data_in(84) xor data_in(87) xor data_in(88) xor data_in(89) xor data_in(91) xor data_in(93) xor data_in(94) xor data_in(96) xor data_in(97) xor data_in(98) xor data_in(100) xor data_in(102) xor data_in(104) xor data_in(105) xor data_in(107) xor data_in(108) xor data_in(113) xor data_in(117) xor data_in(118) xor data_in(121) xor data_in(125) xor data_in(127) xor data_in(128) xor data_in(130) xor data_in(131) xor data_in(133) xor data_in(134) xor data_in(137) xor data_in(138) xor data_in(140) xor data_in(141) xor data_in(143) xor data_in(146) xor data_in(148) xor data_in(149) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(158) xor data_in(161) xor data_in(162) xor data_in(165) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(170) xor data_in(173) xor data_in(174) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(179) xor data_in(181) xor data_in(184) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(191) xor data_in(192) xor data_in(193) xor data_in(194) xor data_in(196) xor data_in(197) xor data_in(199) xor data_in(201) xor data_in(202) xor data_in(204) xor data_in(206) xor data_in(207) xor data_in(210) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(220) xor data_in(221) xor data_in(224) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(232) xor data_in(233) xor data_in(236) xor data_in(237) xor data_in(240) xor data_in(244) xor data_in(245) xor data_in(247) xor data_in(251) xor data_in(252) xor data_in(253) xor data_in(256) xor data_in(258) xor data_in(262) xor data_in(266) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(280) xor data_in(283) xor data_in(286) xor data_in(288) xor data_in(289) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(299) xor data_in(300) xor data_in(305) xor data_in(309) xor data_in(310) xor data_in(311) xor data_in(313) xor data_in(314) xor data_in(317) xor data_in(323) xor data_in(324) xor data_in(325) xor data_in(328) xor data_in(330) xor data_in(332) xor data_in(335) xor data_in(339) xor data_in(340) xor data_in(342) xor data_in(343) xor data_in(344) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(355) xor data_in(356) xor data_in(358) xor data_in(361) xor data_in(365) xor data_in(366) xor data_in(368) xor data_in(371) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(380) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(390) xor data_in(391) xor data_in(395) xor data_in(396) xor data_in(398) xor data_in(399) xor data_in(404) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(417) xor data_in(418) xor data_in(420) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(430) xor data_in(437) xor data_in(439) xor data_in(441) xor data_in(442) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(451) xor data_in(452) xor data_in(453) xor data_in(455) xor data_in(458) xor data_in(460) xor data_in(461) xor data_in(463) xor data_in(465) xor data_in(467) xor data_in(468) xor data_in(470) xor data_in(476) xor data_in(478) xor data_in(482) xor data_in(484) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(495) xor data_in(497) xor data_in(498) xor data_in(502) xor data_in(503) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(509) xor data_in(510) xor data_in(511);
    crc_out(32) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(3) xor crc_in(4) xor crc_in(5) xor crc_in(8) xor crc_in(9) xor crc_in(10) xor crc_in(11) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(22) xor crc_in(23) xor crc_in(24) xor crc_in(25) xor crc_in(26) xor crc_in(28) xor crc_in(29) xor crc_in(30) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(37) xor crc_in(38) xor crc_in(39) xor crc_in(41) xor crc_in(43) xor crc_in(46) xor crc_in(50) xor crc_in(51) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(46) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(65) xor data_in(67) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(73) xor data_in(74) xor data_in(77) xor data_in(80) xor data_in(83) xor data_in(86) xor data_in(87) xor data_in(88) xor data_in(89) xor data_in(90) xor data_in(94) xor data_in(97) xor data_in(98) xor data_in(99) xor data_in(101) xor data_in(102) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(109) xor data_in(110) xor data_in(111) xor data_in(113) xor data_in(118) xor data_in(120) xor data_in(123) xor data_in(124) xor data_in(128) xor data_in(130) xor data_in(131) xor data_in(134) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(140) xor data_in(143) xor data_in(144) xor data_in(146) xor data_in(147) xor data_in(149) xor data_in(151) xor data_in(152) xor data_in(153) xor data_in(157) xor data_in(158) xor data_in(159) xor data_in(160) xor data_in(162) xor data_in(163) xor data_in(164) xor data_in(165) xor data_in(167) xor data_in(169) xor data_in(174) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(184) xor data_in(185) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(192) xor data_in(193) xor data_in(195) xor data_in(198) xor data_in(202) xor data_in(203) xor data_in(204) xor data_in(206) xor data_in(212) xor data_in(214) xor data_in(215) xor data_in(217) xor data_in(218) xor data_in(221) xor data_in(222) xor data_in(223) xor data_in(224) xor data_in(227) xor data_in(232) xor data_in(235) xor data_in(236) xor data_in(238) xor data_in(239) xor data_in(241) xor data_in(242) xor data_in(246) xor data_in(248) xor data_in(253) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(262) xor data_in(264) xor data_in(266) xor data_in(268) xor data_in(269) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(276) xor data_in(278) xor data_in(284) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(293) xor data_in(294) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(304) xor data_in(306) xor data_in(309) xor data_in(310) xor data_in(311) xor data_in(312) xor data_in(313) xor data_in(315) xor data_in(320) xor data_in(323) xor data_in(324) xor data_in(327) xor data_in(329) xor data_in(330) xor data_in(332) xor data_in(334) xor data_in(336) xor data_in(338) xor data_in(339) xor data_in(341) xor data_in(346) xor data_in(348) xor data_in(350) xor data_in(351) xor data_in(353) xor data_in(355) xor data_in(358) xor data_in(359) xor data_in(363) xor data_in(364) xor data_in(366) xor data_in(368) xor data_in(369) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(380) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(387) xor data_in(388) xor data_in(393) xor data_in(395) xor data_in(396) xor data_in(398) xor data_in(399) xor data_in(406) xor data_in(411) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(420) xor data_in(422) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(430) xor data_in(434) xor data_in(435) xor data_in(439) xor data_in(440) xor data_in(443) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(456) xor data_in(460) xor data_in(463) xor data_in(464) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(474) xor data_in(475) xor data_in(478) xor data_in(479) xor data_in(483) xor data_in(484) xor data_in(485) xor data_in(486) xor data_in(489) xor data_in(491) xor data_in(493) xor data_in(505) xor data_in(507) xor data_in(511);
    crc_out(33) <= crc_in(0) xor crc_in(1) xor crc_in(3) xor crc_in(4) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(11) xor crc_in(13) xor crc_in(14) xor crc_in(16) xor crc_in(17) xor crc_in(21) xor crc_in(22) xor crc_in(23) xor crc_in(25) xor crc_in(26) xor crc_in(27) xor crc_in(29) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(38) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(50) xor crc_in(51) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(11) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(25) xor data_in(26) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(50) xor data_in(51) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(63) xor data_in(66) xor data_in(68) xor data_in(69) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(88) xor data_in(89) xor data_in(90) xor data_in(91) xor data_in(92) xor data_in(98) xor data_in(99) xor data_in(100) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(108) xor data_in(112) xor data_in(113) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(125) xor data_in(126) xor data_in(130) xor data_in(131) xor data_in(135) xor data_in(139) xor data_in(140) xor data_in(142) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(151) xor data_in(153) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(159) xor data_in(161) xor data_in(163) xor data_in(167) xor data_in(171) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(184) xor data_in(185) xor data_in(188) xor data_in(189) xor data_in(193) xor data_in(196) xor data_in(197) xor data_in(199) xor data_in(200) xor data_in(203) xor data_in(206) xor data_in(208) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(219) xor data_in(222) xor data_in(226) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(234) xor data_in(235) xor data_in(240) xor data_in(243) xor data_in(245) xor data_in(247) xor data_in(249) xor data_in(252) xor data_in(259) xor data_in(260) xor data_in(262) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(268) xor data_in(270) xor data_in(273) xor data_in(274) xor data_in(276) xor data_in(277) xor data_in(278) xor data_in(279) xor data_in(281) xor data_in(285) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(292) xor data_in(294) xor data_in(297) xor data_in(305) xor data_in(307) xor data_in(309) xor data_in(310) xor data_in(311) xor data_in(312) xor data_in(316) xor data_in(318) xor data_in(320) xor data_in(321) xor data_in(323) xor data_in(324) xor data_in(326) xor data_in(327) xor data_in(328) xor data_in(332) xor data_in(334) xor data_in(335) xor data_in(337) xor data_in(338) xor data_in(342) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(351) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(362) xor data_in(363) xor data_in(365) xor data_in(368) xor data_in(369) xor data_in(370) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(380) xor data_in(381) xor data_in(383) xor data_in(384) xor data_in(387) xor data_in(389) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(398) xor data_in(399) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(413) xor data_in(416) xor data_in(418) xor data_in(420) xor data_in(424) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(430) xor data_in(434) xor data_in(436) xor data_in(438) xor data_in(439) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(444) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(457) xor data_in(459) xor data_in(460) xor data_in(462) xor data_in(463) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(469) xor data_in(474) xor data_in(476) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(480) xor data_in(485) xor data_in(488) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(496) xor data_in(498) xor data_in(499) xor data_in(503) xor data_in(504) xor data_in(505) xor data_in(510);
    crc_out(34) <= crc_in(1) xor crc_in(2) xor crc_in(4) xor crc_in(5) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(10) xor crc_in(12) xor crc_in(14) xor crc_in(15) xor crc_in(17) xor crc_in(18) xor crc_in(22) xor crc_in(23) xor crc_in(24) xor crc_in(26) xor crc_in(27) xor crc_in(28) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(51) xor crc_in(52) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(51) xor data_in(52) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(64) xor data_in(67) xor data_in(69) xor data_in(70) xor data_in(76) xor data_in(77) xor data_in(78) xor data_in(80) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(89) xor data_in(90) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(99) xor data_in(100) xor data_in(101) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(113) xor data_in(114) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(126) xor data_in(127) xor data_in(131) xor data_in(132) xor data_in(136) xor data_in(140) xor data_in(141) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(152) xor data_in(154) xor data_in(156) xor data_in(157) xor data_in(158) xor data_in(160) xor data_in(162) xor data_in(164) xor data_in(168) xor data_in(172) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(185) xor data_in(186) xor data_in(189) xor data_in(190) xor data_in(194) xor data_in(197) xor data_in(198) xor data_in(200) xor data_in(201) xor data_in(204) xor data_in(207) xor data_in(209) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(220) xor data_in(223) xor data_in(227) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(235) xor data_in(236) xor data_in(241) xor data_in(244) xor data_in(246) xor data_in(248) xor data_in(250) xor data_in(253) xor data_in(260) xor data_in(261) xor data_in(263) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(269) xor data_in(271) xor data_in(274) xor data_in(275) xor data_in(277) xor data_in(278) xor data_in(279) xor data_in(280) xor data_in(282) xor data_in(286) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(293) xor data_in(295) xor data_in(298) xor data_in(306) xor data_in(308) xor data_in(310) xor data_in(311) xor data_in(312) xor data_in(313) xor data_in(317) xor data_in(319) xor data_in(321) xor data_in(322) xor data_in(324) xor data_in(325) xor data_in(327) xor data_in(328) xor data_in(329) xor data_in(333) xor data_in(335) xor data_in(336) xor data_in(338) xor data_in(339) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(352) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(363) xor data_in(364) xor data_in(366) xor data_in(369) xor data_in(370) xor data_in(371) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(381) xor data_in(382) xor data_in(384) xor data_in(385) xor data_in(388) xor data_in(390) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(399) xor data_in(400) xor data_in(406) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(414) xor data_in(417) xor data_in(419) xor data_in(421) xor data_in(425) xor data_in(427) xor data_in(428) xor data_in(429) xor data_in(431) xor data_in(435) xor data_in(437) xor data_in(439) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(445) xor data_in(447) xor data_in(448) xor data_in(449) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(458) xor data_in(460) xor data_in(461) xor data_in(463) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(470) xor data_in(475) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(480) xor data_in(481) xor data_in(486) xor data_in(489) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(497) xor data_in(499) xor data_in(500) xor data_in(504) xor data_in(505) xor data_in(506) xor data_in(511);
    crc_out(35) <= crc_in(0) xor crc_in(3) xor crc_in(6) xor crc_in(7) xor crc_in(9) xor crc_in(11) xor crc_in(12) xor crc_in(14) xor crc_in(16) xor crc_in(18) xor crc_in(19) xor crc_in(21) xor crc_in(22) xor crc_in(23) xor crc_in(25) xor crc_in(27) xor crc_in(28) xor crc_in(29) xor crc_in(31) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(37) xor crc_in(40) xor crc_in(42) xor crc_in(44) xor crc_in(46) xor crc_in(50) xor crc_in(54) xor crc_in(55) xor crc_in(60) xor crc_in(61) xor crc_in(63) xor data_in(0) xor data_in(3) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(37) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(46) xor data_in(50) xor data_in(54) xor data_in(55) xor data_in(60) xor data_in(61) xor data_in(63) xor data_in(65) xor data_in(68) xor data_in(69) xor data_in(72) xor data_in(74) xor data_in(76) xor data_in(80) xor data_in(81) xor data_in(84) xor data_in(88) xor data_in(90) xor data_in(91) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(100) xor data_in(101) xor data_in(103) xor data_in(104) xor data_in(106) xor data_in(107) xor data_in(109) xor data_in(111) xor data_in(113) xor data_in(115) xor data_in(119) xor data_in(120) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(128) xor data_in(129) xor data_in(130) xor data_in(133) xor data_in(136) xor data_in(138) xor data_in(139) xor data_in(140) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(156) xor data_in(159) xor data_in(160) xor data_in(161) xor data_in(163) xor data_in(164) xor data_in(166) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(170) xor data_in(171) xor data_in(173) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(180) xor data_in(184) xor data_in(187) xor data_in(191) xor data_in(194) xor data_in(195) xor data_in(197) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(204) xor data_in(206) xor data_in(207) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(215) xor data_in(217) xor data_in(218) xor data_in(221) xor data_in(223) xor data_in(225) xor data_in(226) xor data_in(229) xor data_in(230) xor data_in(235) xor data_in(239) xor data_in(247) xor data_in(249) xor data_in(251) xor data_in(252) xor data_in(258) xor data_in(261) xor data_in(263) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(279) xor data_in(280) xor data_in(283) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(292) xor data_in(294) xor data_in(295) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(300) xor data_in(302) xor data_in(303) xor data_in(304) xor data_in(307) xor data_in(311) xor data_in(312) xor data_in(322) xor data_in(327) xor data_in(328) xor data_in(329) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(336) xor data_in(337) xor data_in(338) xor data_in(343) xor data_in(347) xor data_in(350) xor data_in(352) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(363) xor data_in(365) xor data_in(368) xor data_in(370) xor data_in(371) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(383) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(392) xor data_in(394) xor data_in(396) xor data_in(401) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(424) xor data_in(426) xor data_in(428) xor data_in(431) xor data_in(432) xor data_in(434) xor data_in(435) xor data_in(436) xor data_in(439) xor data_in(440) xor data_in(441) xor data_in(443) xor data_in(444) xor data_in(446) xor data_in(448) xor data_in(450) xor data_in(452) xor data_in(453) xor data_in(455) xor data_in(456) xor data_in(460) xor data_in(463) xor data_in(464) xor data_in(465) xor data_in(467) xor data_in(468) xor data_in(470) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(479) xor data_in(480) xor data_in(481) xor data_in(482) xor data_in(484) xor data_in(486) xor data_in(488) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(494) xor data_in(495) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(503) xor data_in(504) xor data_in(507) xor data_in(508) xor data_in(510);
    crc_out(36) <= crc_in(0) xor crc_in(1) xor crc_in(4) xor crc_in(7) xor crc_in(8) xor crc_in(10) xor crc_in(12) xor crc_in(13) xor crc_in(15) xor crc_in(17) xor crc_in(19) xor crc_in(20) xor crc_in(22) xor crc_in(23) xor crc_in(24) xor crc_in(26) xor crc_in(28) xor crc_in(29) xor crc_in(30) xor crc_in(32) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(38) xor crc_in(41) xor crc_in(43) xor crc_in(45) xor crc_in(47) xor crc_in(51) xor crc_in(55) xor crc_in(56) xor crc_in(61) xor crc_in(62) xor data_in(0) xor data_in(1) xor data_in(4) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(38) xor data_in(41) xor data_in(43) xor data_in(45) xor data_in(47) xor data_in(51) xor data_in(55) xor data_in(56) xor data_in(61) xor data_in(62) xor data_in(64) xor data_in(66) xor data_in(69) xor data_in(70) xor data_in(73) xor data_in(75) xor data_in(77) xor data_in(81) xor data_in(82) xor data_in(85) xor data_in(89) xor data_in(91) xor data_in(92) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(101) xor data_in(102) xor data_in(104) xor data_in(105) xor data_in(107) xor data_in(108) xor data_in(110) xor data_in(112) xor data_in(114) xor data_in(116) xor data_in(120) xor data_in(121) xor data_in(126) xor data_in(127) xor data_in(128) xor data_in(129) xor data_in(130) xor data_in(131) xor data_in(134) xor data_in(137) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(148) xor data_in(149) xor data_in(150) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(157) xor data_in(160) xor data_in(161) xor data_in(162) xor data_in(164) xor data_in(165) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(170) xor data_in(171) xor data_in(172) xor data_in(174) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(181) xor data_in(185) xor data_in(188) xor data_in(192) xor data_in(195) xor data_in(196) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(207) xor data_in(208) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(216) xor data_in(218) xor data_in(219) xor data_in(222) xor data_in(224) xor data_in(226) xor data_in(227) xor data_in(230) xor data_in(231) xor data_in(236) xor data_in(240) xor data_in(248) xor data_in(250) xor data_in(252) xor data_in(253) xor data_in(259) xor data_in(262) xor data_in(264) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(280) xor data_in(281) xor data_in(284) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(293) xor data_in(295) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(301) xor data_in(303) xor data_in(304) xor data_in(305) xor data_in(308) xor data_in(312) xor data_in(313) xor data_in(323) xor data_in(328) xor data_in(329) xor data_in(330) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(337) xor data_in(338) xor data_in(339) xor data_in(344) xor data_in(348) xor data_in(351) xor data_in(353) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(362) xor data_in(364) xor data_in(366) xor data_in(369) xor data_in(371) xor data_in(372) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(384) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(393) xor data_in(395) xor data_in(397) xor data_in(402) xor data_in(406) xor data_in(408) xor data_in(409) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(420) xor data_in(422) xor data_in(423) xor data_in(424) xor data_in(425) xor data_in(427) xor data_in(429) xor data_in(432) xor data_in(433) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(444) xor data_in(445) xor data_in(447) xor data_in(449) xor data_in(451) xor data_in(453) xor data_in(454) xor data_in(456) xor data_in(457) xor data_in(461) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(468) xor data_in(469) xor data_in(471) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(478) xor data_in(480) xor data_in(481) xor data_in(482) xor data_in(483) xor data_in(485) xor data_in(487) xor data_in(489) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(495) xor data_in(496) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(504) xor data_in(505) xor data_in(508) xor data_in(509) xor data_in(511);
    crc_out(37) <= crc_in(0) xor crc_in(1) xor crc_in(7) xor crc_in(9) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(15) xor crc_in(16) xor crc_in(18) xor crc_in(20) xor crc_in(22) xor crc_in(23) xor crc_in(25) xor crc_in(27) xor crc_in(29) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(35) xor crc_in(37) xor crc_in(39) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(47) xor crc_in(48) xor crc_in(50) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(25) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(35) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(50) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(63) xor data_in(65) xor data_in(67) xor data_in(69) xor data_in(72) xor data_in(77) xor data_in(79) xor data_in(80) xor data_in(85) xor data_in(87) xor data_in(90) xor data_in(93) xor data_in(96) xor data_in(97) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(109) xor data_in(110) xor data_in(114) xor data_in(115) xor data_in(117) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(123) xor data_in(124) xor data_in(126) xor data_in(127) xor data_in(128) xor data_in(131) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(139) xor data_in(143) xor data_in(145) xor data_in(147) xor data_in(149) xor data_in(152) xor data_in(153) xor data_in(157) xor data_in(160) xor data_in(161) xor data_in(162) xor data_in(163) xor data_in(164) xor data_in(167) xor data_in(169) xor data_in(172) xor data_in(173) xor data_in(176) xor data_in(181) xor data_in(184) xor data_in(189) xor data_in(190) xor data_in(193) xor data_in(194) xor data_in(196) xor data_in(199) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(207) xor data_in(209) xor data_in(211) xor data_in(213) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(224) xor data_in(226) xor data_in(227) xor data_in(229) xor data_in(230) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(239) xor data_in(241) xor data_in(242) xor data_in(245) xor data_in(249) xor data_in(251) xor data_in(252) xor data_in(253) xor data_in(258) xor data_in(260) xor data_in(262) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(275) xor data_in(276) xor data_in(278) xor data_in(282) xor data_in(285) xor data_in(287) xor data_in(288) xor data_in(290) xor data_in(292) xor data_in(294) xor data_in(295) xor data_in(296) xor data_in(303) xor data_in(305) xor data_in(306) xor data_in(318) xor data_in(320) xor data_in(323) xor data_in(324) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(329) xor data_in(332) xor data_in(335) xor data_in(343) xor data_in(344) xor data_in(346) xor data_in(348) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(360) xor data_in(361) xor data_in(364) xor data_in(365) xor data_in(368) xor data_in(370) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(382) xor data_in(387) xor data_in(389) xor data_in(390) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(400) xor data_in(403) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(410) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(418) xor data_in(425) xor data_in(426) xor data_in(428) xor data_in(429) xor data_in(431) xor data_in(433) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(439) xor data_in(441) xor data_in(443) xor data_in(445) xor data_in(446) xor data_in(448) xor data_in(449) xor data_in(450) xor data_in(453) xor data_in(455) xor data_in(457) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(463) xor data_in(465) xor data_in(467) xor data_in(469) xor data_in(471) xor data_in(472) xor data_in(474) xor data_in(475) xor data_in(476) xor data_in(479) xor data_in(481) xor data_in(482) xor data_in(483) xor data_in(487) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(494) xor data_in(497) xor data_in(498) xor data_in(499) xor data_in(501) xor data_in(502) xor data_in(504) xor data_in(508) xor data_in(509);
    crc_out(38) <= crc_in(1) xor crc_in(2) xor crc_in(8) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(16) xor crc_in(17) xor crc_in(19) xor crc_in(21) xor crc_in(23) xor crc_in(24) xor crc_in(26) xor crc_in(28) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(36) xor crc_in(38) xor crc_in(40) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(47) xor crc_in(48) xor crc_in(49) xor crc_in(51) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor data_in(1) xor data_in(2) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(36) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(49) xor data_in(51) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(64) xor data_in(66) xor data_in(68) xor data_in(70) xor data_in(73) xor data_in(78) xor data_in(80) xor data_in(81) xor data_in(86) xor data_in(88) xor data_in(91) xor data_in(94) xor data_in(97) xor data_in(98) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(110) xor data_in(111) xor data_in(115) xor data_in(116) xor data_in(118) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(124) xor data_in(125) xor data_in(127) xor data_in(128) xor data_in(129) xor data_in(132) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(140) xor data_in(144) xor data_in(146) xor data_in(148) xor data_in(150) xor data_in(153) xor data_in(154) xor data_in(158) xor data_in(161) xor data_in(162) xor data_in(163) xor data_in(164) xor data_in(165) xor data_in(168) xor data_in(170) xor data_in(173) xor data_in(174) xor data_in(177) xor data_in(182) xor data_in(185) xor data_in(190) xor data_in(191) xor data_in(194) xor data_in(195) xor data_in(197) xor data_in(200) xor data_in(202) xor data_in(203) xor data_in(204) xor data_in(206) xor data_in(208) xor data_in(210) xor data_in(212) xor data_in(214) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(225) xor data_in(227) xor data_in(228) xor data_in(230) xor data_in(231) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(240) xor data_in(242) xor data_in(243) xor data_in(246) xor data_in(250) xor data_in(252) xor data_in(253) xor data_in(254) xor data_in(259) xor data_in(261) xor data_in(263) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(273) xor data_in(275) xor data_in(276) xor data_in(277) xor data_in(279) xor data_in(283) xor data_in(286) xor data_in(288) xor data_in(289) xor data_in(291) xor data_in(293) xor data_in(295) xor data_in(296) xor data_in(297) xor data_in(304) xor data_in(306) xor data_in(307) xor data_in(319) xor data_in(321) xor data_in(324) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(328) xor data_in(330) xor data_in(333) xor data_in(336) xor data_in(344) xor data_in(345) xor data_in(347) xor data_in(349) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(361) xor data_in(362) xor data_in(365) xor data_in(366) xor data_in(369) xor data_in(371) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(383) xor data_in(388) xor data_in(390) xor data_in(391) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(398) xor data_in(401) xor data_in(404) xor data_in(406) xor data_in(408) xor data_in(409) xor data_in(411) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(419) xor data_in(426) xor data_in(427) xor data_in(429) xor data_in(430) xor data_in(432) xor data_in(434) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(440) xor data_in(442) xor data_in(444) xor data_in(446) xor data_in(447) xor data_in(449) xor data_in(450) xor data_in(451) xor data_in(454) xor data_in(456) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(464) xor data_in(466) xor data_in(468) xor data_in(470) xor data_in(472) xor data_in(473) xor data_in(475) xor data_in(476) xor data_in(477) xor data_in(480) xor data_in(482) xor data_in(483) xor data_in(484) xor data_in(488) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(495) xor data_in(498) xor data_in(499) xor data_in(500) xor data_in(502) xor data_in(503) xor data_in(505) xor data_in(509) xor data_in(510);
    crc_out(39) <= crc_in(0) xor crc_in(2) xor crc_in(3) xor crc_in(9) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(17) xor crc_in(18) xor crc_in(20) xor crc_in(22) xor crc_in(24) xor crc_in(25) xor crc_in(27) xor crc_in(29) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(37) xor crc_in(39) xor crc_in(41) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(47) xor crc_in(48) xor crc_in(49) xor crc_in(50) xor crc_in(52) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor data_in(0) xor data_in(2) xor data_in(3) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(22) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(52) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(65) xor data_in(67) xor data_in(69) xor data_in(71) xor data_in(74) xor data_in(79) xor data_in(81) xor data_in(82) xor data_in(87) xor data_in(89) xor data_in(92) xor data_in(95) xor data_in(98) xor data_in(99) xor data_in(106) xor data_in(107) xor data_in(108) xor data_in(111) xor data_in(112) xor data_in(116) xor data_in(117) xor data_in(119) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(125) xor data_in(126) xor data_in(128) xor data_in(129) xor data_in(130) xor data_in(133) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(141) xor data_in(145) xor data_in(147) xor data_in(149) xor data_in(151) xor data_in(154) xor data_in(155) xor data_in(159) xor data_in(162) xor data_in(163) xor data_in(164) xor data_in(165) xor data_in(166) xor data_in(169) xor data_in(171) xor data_in(174) xor data_in(175) xor data_in(178) xor data_in(183) xor data_in(186) xor data_in(191) xor data_in(192) xor data_in(195) xor data_in(196) xor data_in(198) xor data_in(201) xor data_in(203) xor data_in(204) xor data_in(205) xor data_in(207) xor data_in(209) xor data_in(211) xor data_in(213) xor data_in(215) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(226) xor data_in(228) xor data_in(229) xor data_in(231) xor data_in(232) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(241) xor data_in(243) xor data_in(244) xor data_in(247) xor data_in(251) xor data_in(253) xor data_in(254) xor data_in(255) xor data_in(260) xor data_in(262) xor data_in(264) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(274) xor data_in(276) xor data_in(277) xor data_in(278) xor data_in(280) xor data_in(284) xor data_in(287) xor data_in(289) xor data_in(290) xor data_in(292) xor data_in(294) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(305) xor data_in(307) xor data_in(308) xor data_in(320) xor data_in(322) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(328) xor data_in(329) xor data_in(331) xor data_in(334) xor data_in(337) xor data_in(345) xor data_in(346) xor data_in(348) xor data_in(350) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(359) xor data_in(360) xor data_in(362) xor data_in(363) xor data_in(366) xor data_in(367) xor data_in(370) xor data_in(372) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(380) xor data_in(384) xor data_in(389) xor data_in(391) xor data_in(392) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(398) xor data_in(399) xor data_in(402) xor data_in(405) xor data_in(407) xor data_in(409) xor data_in(410) xor data_in(412) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(420) xor data_in(427) xor data_in(428) xor data_in(430) xor data_in(431) xor data_in(433) xor data_in(435) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(441) xor data_in(443) xor data_in(445) xor data_in(447) xor data_in(448) xor data_in(450) xor data_in(451) xor data_in(452) xor data_in(455) xor data_in(457) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(463) xor data_in(465) xor data_in(467) xor data_in(469) xor data_in(471) xor data_in(473) xor data_in(474) xor data_in(476) xor data_in(477) xor data_in(478) xor data_in(481) xor data_in(483) xor data_in(484) xor data_in(485) xor data_in(489) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(496) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(503) xor data_in(504) xor data_in(506) xor data_in(510) xor data_in(511);
    crc_out(40) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(3) xor crc_in(4) xor crc_in(5) xor crc_in(7) xor crc_in(8) xor crc_in(18) xor crc_in(19) xor crc_in(22) xor crc_in(23) xor crc_in(24) xor crc_in(25) xor crc_in(26) xor crc_in(28) xor crc_in(30) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(38) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(46) xor crc_in(48) xor crc_in(49) xor crc_in(51) xor crc_in(52) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(60) xor crc_in(61) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(18) xor data_in(19) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(30) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(38) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(48) xor data_in(49) xor data_in(51) xor data_in(52) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(60) xor data_in(61) xor data_in(66) xor data_in(68) xor data_in(69) xor data_in(71) xor data_in(74) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(88) xor data_in(90) xor data_in(92) xor data_in(93) xor data_in(95) xor data_in(96) xor data_in(99) xor data_in(100) xor data_in(102) xor data_in(103) xor data_in(104) xor data_in(107) xor data_in(109) xor data_in(110) xor data_in(111) xor data_in(112) xor data_in(114) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(127) xor data_in(131) xor data_in(132) xor data_in(134) xor data_in(136) xor data_in(137) xor data_in(141) xor data_in(143) xor data_in(148) xor data_in(151) xor data_in(154) xor data_in(157) xor data_in(158) xor data_in(163) xor data_in(168) xor data_in(171) xor data_in(172) xor data_in(177) xor data_in(178) xor data_in(181) xor data_in(182) xor data_in(186) xor data_in(187) xor data_in(190) xor data_in(192) xor data_in(193) xor data_in(194) xor data_in(196) xor data_in(199) xor data_in(200) xor data_in(202) xor data_in(207) xor data_in(210) xor data_in(211) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(224) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(231) xor data_in(234) xor data_in(235) xor data_in(238) xor data_in(244) xor data_in(248) xor data_in(255) xor data_in(256) xor data_in(258) xor data_in(261) xor data_in(262) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(276) xor data_in(277) xor data_in(279) xor data_in(285) xor data_in(287) xor data_in(290) xor data_in(293) xor data_in(300) xor data_in(302) xor data_in(303) xor data_in(304) xor data_in(306) xor data_in(308) xor data_in(313) xor data_in(314) xor data_in(318) xor data_in(320) xor data_in(321) xor data_in(325) xor data_in(328) xor data_in(329) xor data_in(331) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(339) xor data_in(340) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(347) xor data_in(348) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(355) xor data_in(359) xor data_in(360) xor data_in(361) xor data_in(362) xor data_in(371) xor data_in(372) xor data_in(378) xor data_in(381) xor data_in(382) xor data_in(387) xor data_in(388) xor data_in(390) xor data_in(391) xor data_in(396) xor data_in(399) xor data_in(403) xor data_in(405) xor data_in(406) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(416) xor data_in(418) xor data_in(420) xor data_in(423) xor data_in(424) xor data_in(428) xor data_in(430) xor data_in(432) xor data_in(435) xor data_in(436) xor data_in(440) xor data_in(444) xor data_in(446) xor data_in(448) xor data_in(451) xor data_in(454) xor data_in(456) xor data_in(458) xor data_in(459) xor data_in(464) xor data_in(468) xor data_in(471) xor data_in(472) xor data_in(479) xor data_in(482) xor data_in(485) xor data_in(487) xor data_in(488) xor data_in(490) xor data_in(491) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(497) xor data_in(498) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(503) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(510) xor data_in(511);
    crc_out(41) <= crc_in(0) xor crc_in(1) xor crc_in(3) xor crc_in(4) xor crc_in(6) xor crc_in(7) xor crc_in(9) xor crc_in(10) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(19) xor crc_in(20) xor crc_in(21) xor crc_in(22) xor crc_in(23) xor crc_in(25) xor crc_in(26) xor crc_in(27) xor crc_in(29) xor crc_in(31) xor crc_in(32) xor crc_in(34) xor crc_in(35) xor crc_in(39) xor crc_in(42) xor crc_in(44) xor crc_in(49) xor crc_in(54) xor crc_in(56) xor crc_in(57) xor crc_in(59) xor crc_in(61) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(25) xor data_in(26) xor data_in(27) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(39) xor data_in(42) xor data_in(44) xor data_in(49) xor data_in(54) xor data_in(56) xor data_in(57) xor data_in(59) xor data_in(61) xor data_in(67) xor data_in(71) xor data_in(74) xor data_in(75) xor data_in(82) xor data_in(83) xor data_in(85) xor data_in(88) xor data_in(89) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(97) xor data_in(100) xor data_in(101) xor data_in(102) xor data_in(105) xor data_in(112) xor data_in(114) xor data_in(115) xor data_in(118) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(126) xor data_in(128) xor data_in(129) xor data_in(130) xor data_in(133) xor data_in(135) xor data_in(136) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(143) xor data_in(144) xor data_in(146) xor data_in(149) xor data_in(150) xor data_in(151) xor data_in(154) xor data_in(156) xor data_in(157) xor data_in(159) xor data_in(160) xor data_in(165) xor data_in(166) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(170) xor data_in(171) xor data_in(172) xor data_in(173) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(181) xor data_in(183) xor data_in(184) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(190) xor data_in(191) xor data_in(193) xor data_in(195) xor data_in(201) xor data_in(203) xor data_in(204) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(214) xor data_in(216) xor data_in(218) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(224) xor data_in(227) xor data_in(230) xor data_in(231) xor data_in(233) xor data_in(234) xor data_in(237) xor data_in(242) xor data_in(249) xor data_in(252) xor data_in(254) xor data_in(256) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(264) xor data_in(265) xor data_in(268) xor data_in(269) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(276) xor data_in(277) xor data_in(280) xor data_in(281) xor data_in(286) xor data_in(287) xor data_in(294) xor data_in(295) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(305) xor data_in(307) xor data_in(313) xor data_in(315) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(325) xor data_in(327) xor data_in(329) xor data_in(331) xor data_in(333) xor data_in(335) xor data_in(336) xor data_in(338) xor data_in(339) xor data_in(341) xor data_in(343) xor data_in(354) xor data_in(355) xor data_in(357) xor data_in(358) xor data_in(360) xor data_in(361) xor data_in(364) xor data_in(367) xor data_in(368) xor data_in(380) xor data_in(383) xor data_in(385) xor data_in(387) xor data_in(389) xor data_in(393) xor data_in(395) xor data_in(398) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(411) xor data_in(416) xor data_in(420) xor data_in(423) xor data_in(425) xor data_in(430) xor data_in(433) xor data_in(434) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(441) xor data_in(442) xor data_in(445) xor data_in(447) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(457) xor data_in(461) xor data_in(462) xor data_in(463) xor data_in(465) xor data_in(466) xor data_in(469) xor data_in(470) xor data_in(471) xor data_in(472) xor data_in(473) xor data_in(474) xor data_in(475) xor data_in(477) xor data_in(478) xor data_in(480) xor data_in(483) xor data_in(484) xor data_in(487) xor data_in(489) xor data_in(492) xor data_in(493) xor data_in(495) xor data_in(497) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(509) xor data_in(510) xor data_in(511);
    crc_out(42) <= crc_in(0) xor crc_in(1) xor crc_in(4) xor crc_in(11) xor crc_in(12) xor crc_in(16) xor crc_in(20) xor crc_in(23) xor crc_in(26) xor crc_in(27) xor crc_in(28) xor crc_in(30) xor crc_in(33) xor crc_in(35) xor crc_in(40) xor crc_in(41) xor crc_in(47) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(57) xor crc_in(59) xor crc_in(60) xor data_in(0) xor data_in(1) xor data_in(4) xor data_in(11) xor data_in(12) xor data_in(16) xor data_in(20) xor data_in(23) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(33) xor data_in(35) xor data_in(40) xor data_in(41) xor data_in(47) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(57) xor data_in(59) xor data_in(60) xor data_in(68) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(74) xor data_in(75) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(82) xor data_in(84) xor data_in(85) xor data_in(87) xor data_in(89) xor data_in(90) xor data_in(93) xor data_in(94) xor data_in(96) xor data_in(97) xor data_in(98) xor data_in(101) xor data_in(104) xor data_in(106) xor data_in(108) xor data_in(110) xor data_in(111) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(120) xor data_in(122) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(131) xor data_in(132) xor data_in(134) xor data_in(138) xor data_in(139) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(147) xor data_in(154) xor data_in(156) xor data_in(161) xor data_in(164) xor data_in(165) xor data_in(169) xor data_in(172) xor data_in(173) xor data_in(174) xor data_in(175) xor data_in(179) xor data_in(181) xor data_in(185) xor data_in(186) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(190) xor data_in(191) xor data_in(192) xor data_in(196) xor data_in(197) xor data_in(200) xor data_in(202) xor data_in(211) xor data_in(212) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(221) xor data_in(222) xor data_in(224) xor data_in(226) xor data_in(229) xor data_in(230) xor data_in(233) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(239) xor data_in(242) xor data_in(243) xor data_in(245) xor data_in(250) xor data_in(252) xor data_in(253) xor data_in(254) xor data_in(255) xor data_in(257) xor data_in(259) xor data_in(260) xor data_in(262) xor data_in(263) xor data_in(264) xor data_in(265) xor data_in(267) xor data_in(268) xor data_in(270) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(275) xor data_in(276) xor data_in(277) xor data_in(282) xor data_in(291) xor data_in(296) xor data_in(297) xor data_in(301) xor data_in(304) xor data_in(306) xor data_in(308) xor data_in(309) xor data_in(313) xor data_in(316) xor data_in(318) xor data_in(319) xor data_in(321) xor data_in(322) xor data_in(324) xor data_in(325) xor data_in(327) xor data_in(328) xor data_in(331) xor data_in(333) xor data_in(336) xor data_in(337) xor data_in(338) xor data_in(342) xor data_in(343) xor data_in(345) xor data_in(346) xor data_in(348) xor data_in(349) xor data_in(352) xor data_in(353) xor data_in(357) xor data_in(359) xor data_in(361) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(367) xor data_in(369) xor data_in(372) xor data_in(373) xor data_in(379) xor data_in(380) xor data_in(381) xor data_in(382) xor data_in(384) xor data_in(385) xor data_in(386) xor data_in(387) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(406) xor data_in(407) xor data_in(410) xor data_in(411) xor data_in(413) xor data_in(416) xor data_in(419) xor data_in(420) xor data_in(423) xor data_in(426) xor data_in(429) xor data_in(430) xor data_in(436) xor data_in(437) xor data_in(440) xor data_in(443) xor data_in(446) xor data_in(448) xor data_in(449) xor data_in(452) xor data_in(453) xor data_in(455) xor data_in(456) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(464) xor data_in(467) xor data_in(472) xor data_in(473) xor data_in(476) xor data_in(477) xor data_in(479) xor data_in(481) xor data_in(485) xor data_in(486) xor data_in(487) xor data_in(490) xor data_in(491) xor data_in(494) xor data_in(499) xor data_in(501) xor data_in(502) xor data_in(504) xor data_in(505) xor data_in(507) xor data_in(511);
    crc_out(43) <= crc_in(0) xor crc_in(1) xor crc_in(7) xor crc_in(8) xor crc_in(10) xor crc_in(14) xor crc_in(15) xor crc_in(17) xor crc_in(22) xor crc_in(27) xor crc_in(28) xor crc_in(29) xor crc_in(31) xor crc_in(32) xor crc_in(34) xor crc_in(42) xor crc_in(43) xor crc_in(45) xor crc_in(47) xor crc_in(48) xor crc_in(50) xor crc_in(52) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor data_in(0) xor data_in(1) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(22) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(34) xor data_in(42) xor data_in(43) xor data_in(45) xor data_in(47) xor data_in(48) xor data_in(50) xor data_in(52) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(74) xor data_in(75) xor data_in(77) xor data_in(81) xor data_in(82) xor data_in(87) xor data_in(88) xor data_in(90) xor data_in(91) xor data_in(92) xor data_in(94) xor data_in(97) xor data_in(98) xor data_in(99) xor data_in(103) xor data_in(104) xor data_in(105) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(112) xor data_in(113) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(124) xor data_in(127) xor data_in(128) xor data_in(129) xor data_in(130) xor data_in(133) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(141) xor data_in(142) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(147) xor data_in(148) xor data_in(150) xor data_in(151) xor data_in(152) xor data_in(154) xor data_in(156) xor data_in(158) xor data_in(160) xor data_in(162) xor data_in(164) xor data_in(167) xor data_in(168) xor data_in(171) xor data_in(173) xor data_in(174) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(184) xor data_in(187) xor data_in(188) xor data_in(189) xor data_in(191) xor data_in(192) xor data_in(193) xor data_in(194) xor data_in(198) xor data_in(200) xor data_in(201) xor data_in(203) xor data_in(204) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(208) xor data_in(211) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(217) xor data_in(219) xor data_in(220) xor data_in(222) xor data_in(224) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(232) xor data_in(233) xor data_in(235) xor data_in(236) xor data_in(238) xor data_in(240) xor data_in(242) xor data_in(243) xor data_in(244) xor data_in(245) xor data_in(246) xor data_in(251) xor data_in(252) xor data_in(253) xor data_in(255) xor data_in(256) xor data_in(260) xor data_in(261) xor data_in(262) xor data_in(265) xor data_in(267) xor data_in(271) xor data_in(273) xor data_in(274) xor data_in(277) xor data_in(281) xor data_in(283) xor data_in(287) xor data_in(288) xor data_in(291) xor data_in(292) xor data_in(295) xor data_in(299) xor data_in(300) xor data_in(303) xor data_in(304) xor data_in(305) xor data_in(307) xor data_in(310) xor data_in(313) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(322) xor data_in(327) xor data_in(328) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(333) xor data_in(337) xor data_in(340) xor data_in(345) xor data_in(347) xor data_in(348) xor data_in(350) xor data_in(352) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(360) xor data_in(363) xor data_in(365) xor data_in(366) xor data_in(367) xor data_in(370) xor data_in(372) xor data_in(374) xor data_in(379) xor data_in(381) xor data_in(383) xor data_in(386) xor data_in(394) xor data_in(396) xor data_in(399) xor data_in(401) xor data_in(405) xor data_in(407) xor data_in(409) xor data_in(411) xor data_in(413) xor data_in(414) xor data_in(416) xor data_in(419) xor data_in(423) xor data_in(427) xor data_in(429) xor data_in(434) xor data_in(435) xor data_in(437) xor data_in(439) xor data_in(441) xor data_in(442) xor data_in(444) xor data_in(447) xor data_in(450) xor data_in(452) xor data_in(456) xor data_in(457) xor data_in(463) xor data_in(465) xor data_in(466) xor data_in(468) xor data_in(470) xor data_in(471) xor data_in(473) xor data_in(475) xor data_in(480) xor data_in(482) xor data_in(484) xor data_in(492) xor data_in(493) xor data_in(495) xor data_in(496) xor data_in(498) xor data_in(499) xor data_in(500) xor data_in(502) xor data_in(504) xor data_in(510);
    crc_out(44) <= crc_in(1) xor crc_in(2) xor crc_in(8) xor crc_in(9) xor crc_in(11) xor crc_in(15) xor crc_in(16) xor crc_in(18) xor crc_in(23) xor crc_in(28) xor crc_in(29) xor crc_in(30) xor crc_in(32) xor crc_in(33) xor crc_in(35) xor crc_in(43) xor crc_in(44) xor crc_in(46) xor crc_in(48) xor crc_in(49) xor crc_in(51) xor crc_in(53) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(1) xor data_in(2) xor data_in(8) xor data_in(9) xor data_in(11) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(23) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(33) xor data_in(35) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(48) xor data_in(49) xor data_in(51) xor data_in(53) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(75) xor data_in(76) xor data_in(78) xor data_in(82) xor data_in(83) xor data_in(88) xor data_in(89) xor data_in(91) xor data_in(92) xor data_in(93) xor data_in(95) xor data_in(98) xor data_in(99) xor data_in(100) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(111) xor data_in(113) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(125) xor data_in(128) xor data_in(129) xor data_in(130) xor data_in(131) xor data_in(134) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(142) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(146) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(157) xor data_in(159) xor data_in(161) xor data_in(163) xor data_in(165) xor data_in(168) xor data_in(169) xor data_in(172) xor data_in(174) xor data_in(175) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(185) xor data_in(188) xor data_in(189) xor data_in(190) xor data_in(192) xor data_in(193) xor data_in(194) xor data_in(195) xor data_in(199) xor data_in(201) xor data_in(202) xor data_in(204) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(208) xor data_in(209) xor data_in(212) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(218) xor data_in(220) xor data_in(221) xor data_in(223) xor data_in(225) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(233) xor data_in(234) xor data_in(236) xor data_in(237) xor data_in(239) xor data_in(241) xor data_in(243) xor data_in(244) xor data_in(245) xor data_in(246) xor data_in(247) xor data_in(252) xor data_in(253) xor data_in(254) xor data_in(256) xor data_in(257) xor data_in(261) xor data_in(262) xor data_in(263) xor data_in(266) xor data_in(268) xor data_in(272) xor data_in(274) xor data_in(275) xor data_in(278) xor data_in(282) xor data_in(284) xor data_in(288) xor data_in(289) xor data_in(292) xor data_in(293) xor data_in(296) xor data_in(300) xor data_in(301) xor data_in(304) xor data_in(305) xor data_in(306) xor data_in(308) xor data_in(311) xor data_in(314) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(323) xor data_in(328) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(334) xor data_in(338) xor data_in(341) xor data_in(346) xor data_in(348) xor data_in(349) xor data_in(351) xor data_in(353) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(358) xor data_in(361) xor data_in(364) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(371) xor data_in(373) xor data_in(375) xor data_in(380) xor data_in(382) xor data_in(384) xor data_in(387) xor data_in(395) xor data_in(397) xor data_in(400) xor data_in(402) xor data_in(406) xor data_in(408) xor data_in(410) xor data_in(412) xor data_in(414) xor data_in(415) xor data_in(417) xor data_in(420) xor data_in(424) xor data_in(428) xor data_in(430) xor data_in(435) xor data_in(436) xor data_in(438) xor data_in(440) xor data_in(442) xor data_in(443) xor data_in(445) xor data_in(448) xor data_in(451) xor data_in(453) xor data_in(457) xor data_in(458) xor data_in(464) xor data_in(466) xor data_in(467) xor data_in(469) xor data_in(471) xor data_in(472) xor data_in(474) xor data_in(476) xor data_in(481) xor data_in(483) xor data_in(485) xor data_in(493) xor data_in(494) xor data_in(496) xor data_in(497) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(503) xor data_in(505) xor data_in(511);
    crc_out(45) <= crc_in(0) xor crc_in(3) xor crc_in(5) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(17) xor crc_in(19) xor crc_in(21) xor crc_in(22) xor crc_in(29) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(41) xor crc_in(43) xor crc_in(44) xor crc_in(49) xor crc_in(53) xor crc_in(55) xor crc_in(58) xor crc_in(59) xor crc_in(61) xor crc_in(63) xor data_in(0) xor data_in(3) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(49) xor data_in(53) xor data_in(55) xor data_in(58) xor data_in(59) xor data_in(61) xor data_in(63) xor data_in(64) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(74) xor data_in(78) xor data_in(80) xor data_in(82) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(89) xor data_in(90) xor data_in(93) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(99) xor data_in(100) xor data_in(101) xor data_in(102) xor data_in(103) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(112) xor data_in(113) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(120) xor data_in(121) xor data_in(131) xor data_in(135) xor data_in(136) xor data_in(141) xor data_in(142) xor data_in(144) xor data_in(145) xor data_in(147) xor data_in(149) xor data_in(151) xor data_in(153) xor data_in(155) xor data_in(157) xor data_in(162) xor data_in(165) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(171) xor data_in(173) xor data_in(177) xor data_in(178) xor data_in(180) xor data_in(183) xor data_in(184) xor data_in(189) xor data_in(191) xor data_in(193) xor data_in(195) xor data_in(196) xor data_in(197) xor data_in(202) xor data_in(203) xor data_in(204) xor data_in(209) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(221) xor data_in(222) xor data_in(223) xor data_in(225) xor data_in(232) xor data_in(233) xor data_in(236) xor data_in(238) xor data_in(239) xor data_in(240) xor data_in(244) xor data_in(246) xor data_in(247) xor data_in(248) xor data_in(252) xor data_in(253) xor data_in(255) xor data_in(257) xor data_in(266) xor data_in(268) xor data_in(273) xor data_in(278) xor data_in(279) xor data_in(281) xor data_in(283) xor data_in(285) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(293) xor data_in(294) xor data_in(295) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(303) xor data_in(304) xor data_in(305) xor data_in(306) xor data_in(307) xor data_in(312) xor data_in(313) xor data_in(314) xor data_in(315) xor data_in(318) xor data_in(319) xor data_in(321) xor data_in(323) xor data_in(324) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(329) xor data_in(334) xor data_in(335) xor data_in(338) xor data_in(340) xor data_in(342) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(350) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(359) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(369) xor data_in(373) xor data_in(374) xor data_in(376) xor data_in(379) xor data_in(380) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(387) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(400) xor data_in(401) xor data_in(403) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(411) xor data_in(412) xor data_in(415) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(420) xor data_in(423) xor data_in(424) xor data_in(425) xor data_in(430) xor data_in(434) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(446) xor data_in(453) xor data_in(458) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(463) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(471) xor data_in(472) xor data_in(473) xor data_in(474) xor data_in(478) xor data_in(482) xor data_in(487) xor data_in(488) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(497) xor data_in(499) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(503) xor data_in(505) xor data_in(508) xor data_in(510);
    crc_out(46) <= crc_in(0) xor crc_in(1) xor crc_in(4) xor crc_in(6) xor crc_in(8) xor crc_in(9) xor crc_in(10) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(17) xor crc_in(18) xor crc_in(20) xor crc_in(22) xor crc_in(23) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(42) xor crc_in(44) xor crc_in(45) xor crc_in(50) xor crc_in(54) xor crc_in(56) xor crc_in(59) xor crc_in(60) xor crc_in(62) xor data_in(0) xor data_in(1) xor data_in(4) xor data_in(6) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(42) xor data_in(44) xor data_in(45) xor data_in(50) xor data_in(54) xor data_in(56) xor data_in(59) xor data_in(60) xor data_in(62) xor data_in(64) xor data_in(65) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(75) xor data_in(79) xor data_in(81) xor data_in(83) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(88) xor data_in(90) xor data_in(91) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(97) xor data_in(100) xor data_in(101) xor data_in(102) xor data_in(103) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(113) xor data_in(114) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(121) xor data_in(122) xor data_in(132) xor data_in(136) xor data_in(137) xor data_in(142) xor data_in(143) xor data_in(145) xor data_in(146) xor data_in(148) xor data_in(150) xor data_in(152) xor data_in(154) xor data_in(156) xor data_in(158) xor data_in(163) xor data_in(166) xor data_in(168) xor data_in(169) xor data_in(170) xor data_in(172) xor data_in(174) xor data_in(178) xor data_in(179) xor data_in(181) xor data_in(184) xor data_in(185) xor data_in(190) xor data_in(192) xor data_in(194) xor data_in(196) xor data_in(197) xor data_in(198) xor data_in(203) xor data_in(204) xor data_in(205) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(222) xor data_in(223) xor data_in(224) xor data_in(226) xor data_in(233) xor data_in(234) xor data_in(237) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(245) xor data_in(247) xor data_in(248) xor data_in(249) xor data_in(253) xor data_in(254) xor data_in(256) xor data_in(258) xor data_in(267) xor data_in(269) xor data_in(274) xor data_in(279) xor data_in(280) xor data_in(282) xor data_in(284) xor data_in(286) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(294) xor data_in(295) xor data_in(296) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(304) xor data_in(305) xor data_in(306) xor data_in(307) xor data_in(308) xor data_in(313) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(319) xor data_in(320) xor data_in(322) xor data_in(324) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(328) xor data_in(330) xor data_in(335) xor data_in(336) xor data_in(339) xor data_in(341) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(351) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(360) xor data_in(364) xor data_in(365) xor data_in(366) xor data_in(370) xor data_in(374) xor data_in(375) xor data_in(377) xor data_in(380) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(388) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(396) xor data_in(397) xor data_in(398) xor data_in(401) xor data_in(402) xor data_in(404) xor data_in(406) xor data_in(408) xor data_in(409) xor data_in(412) xor data_in(413) xor data_in(416) xor data_in(418) xor data_in(419) xor data_in(420) xor data_in(421) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(431) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(447) xor data_in(454) xor data_in(459) xor data_in(461) xor data_in(462) xor data_in(463) xor data_in(464) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(472) xor data_in(473) xor data_in(474) xor data_in(475) xor data_in(479) xor data_in(483) xor data_in(488) xor data_in(489) xor data_in(492) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(497) xor data_in(498) xor data_in(500) xor data_in(501) xor data_in(502) xor data_in(503) xor data_in(504) xor data_in(506) xor data_in(509) xor data_in(511);
    crc_out(47) <= crc_in(0) xor crc_in(1) xor crc_in(8) xor crc_in(9) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(16) xor crc_in(17) xor crc_in(18) xor crc_in(19) xor crc_in(22) xor crc_in(23) xor crc_in(31) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(41) xor crc_in(46) xor crc_in(47) xor crc_in(50) xor crc_in(51) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(57) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(8) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(22) xor data_in(23) xor data_in(31) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(41) xor data_in(46) xor data_in(47) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(65) xor data_in(66) xor data_in(69) xor data_in(70) xor data_in(73) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(88) xor data_in(89) xor data_in(91) xor data_in(96) xor data_in(97) xor data_in(98) xor data_in(101) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(109) xor data_in(113) xor data_in(115) xor data_in(117) xor data_in(118) xor data_in(124) xor data_in(126) xor data_in(129) xor data_in(130) xor data_in(132) xor data_in(133) xor data_in(136) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(142) xor data_in(144) xor data_in(147) xor data_in(149) xor data_in(150) xor data_in(152) xor data_in(153) xor data_in(154) xor data_in(156) xor data_in(158) xor data_in(159) xor data_in(160) xor data_in(165) xor data_in(166) xor data_in(168) xor data_in(169) xor data_in(173) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(180) xor data_in(181) xor data_in(184) xor data_in(185) xor data_in(190) xor data_in(191) xor data_in(193) xor data_in(194) xor data_in(195) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(207) xor data_in(208) xor data_in(213) xor data_in(215) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(245) xor data_in(246) xor data_in(248) xor data_in(249) xor data_in(250) xor data_in(252) xor data_in(255) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(262) xor data_in(263) xor data_in(264) xor data_in(266) xor data_in(267) xor data_in(269) xor data_in(270) xor data_in(276) xor data_in(278) xor data_in(280) xor data_in(283) xor data_in(285) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(292) xor data_in(293) xor data_in(296) xor data_in(298) xor data_in(299) xor data_in(301) xor data_in(304) xor data_in(305) xor data_in(306) xor data_in(307) xor data_in(308) xor data_in(313) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(321) xor data_in(328) xor data_in(329) xor data_in(330) xor data_in(332) xor data_in(333) xor data_in(334) xor data_in(336) xor data_in(337) xor data_in(338) xor data_in(339) xor data_in(342) xor data_in(343) xor data_in(347) xor data_in(350) xor data_in(353) xor data_in(358) xor data_in(361) xor data_in(362) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(366) xor data_in(368) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(375) xor data_in(376) xor data_in(378) xor data_in(379) xor data_in(380) xor data_in(381) xor data_in(383) xor data_in(384) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(391) xor data_in(392) xor data_in(394) xor data_in(399) xor data_in(400) xor data_in(402) xor data_in(403) xor data_in(407) xor data_in(408) xor data_in(410) xor data_in(412) xor data_in(414) xor data_in(416) xor data_in(422) xor data_in(423) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(429) xor data_in(430) xor data_in(431) xor data_in(432) xor data_in(434) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(440) xor data_in(442) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(448) xor data_in(449) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(459) xor data_in(461) xor data_in(464) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(471) xor data_in(473) xor data_in(476) xor data_in(477) xor data_in(478) xor data_in(480) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(495) xor data_in(497) xor data_in(501) xor data_in(502) xor data_in(506) xor data_in(507) xor data_in(508);
    crc_out(48) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(9) xor crc_in(10) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(17) xor crc_in(18) xor crc_in(19) xor crc_in(20) xor crc_in(23) xor crc_in(24) xor crc_in(32) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(42) xor crc_in(47) xor crc_in(48) xor crc_in(51) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(58) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(23) xor data_in(24) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(42) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(64) xor data_in(66) xor data_in(67) xor data_in(70) xor data_in(71) xor data_in(74) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(89) xor data_in(90) xor data_in(92) xor data_in(97) xor data_in(98) xor data_in(99) xor data_in(102) xor data_in(106) xor data_in(107) xor data_in(108) xor data_in(110) xor data_in(114) xor data_in(116) xor data_in(118) xor data_in(119) xor data_in(125) xor data_in(127) xor data_in(130) xor data_in(131) xor data_in(133) xor data_in(134) xor data_in(137) xor data_in(140) xor data_in(141) xor data_in(142) xor data_in(143) xor data_in(145) xor data_in(148) xor data_in(150) xor data_in(151) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(157) xor data_in(159) xor data_in(160) xor data_in(161) xor data_in(166) xor data_in(167) xor data_in(169) xor data_in(170) xor data_in(174) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(181) xor data_in(182) xor data_in(185) xor data_in(186) xor data_in(191) xor data_in(192) xor data_in(194) xor data_in(195) xor data_in(196) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(208) xor data_in(209) xor data_in(214) xor data_in(216) xor data_in(218) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(237) xor data_in(238) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(242) xor data_in(246) xor data_in(247) xor data_in(249) xor data_in(250) xor data_in(251) xor data_in(253) xor data_in(256) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(263) xor data_in(264) xor data_in(265) xor data_in(267) xor data_in(268) xor data_in(270) xor data_in(271) xor data_in(277) xor data_in(279) xor data_in(281) xor data_in(284) xor data_in(286) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(293) xor data_in(294) xor data_in(297) xor data_in(299) xor data_in(300) xor data_in(302) xor data_in(305) xor data_in(306) xor data_in(307) xor data_in(308) xor data_in(309) xor data_in(314) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(322) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(337) xor data_in(338) xor data_in(339) xor data_in(340) xor data_in(343) xor data_in(344) xor data_in(348) xor data_in(351) xor data_in(354) xor data_in(359) xor data_in(362) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(366) xor data_in(367) xor data_in(369) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(376) xor data_in(377) xor data_in(379) xor data_in(380) xor data_in(381) xor data_in(382) xor data_in(384) xor data_in(385) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(392) xor data_in(393) xor data_in(395) xor data_in(400) xor data_in(401) xor data_in(403) xor data_in(404) xor data_in(408) xor data_in(409) xor data_in(411) xor data_in(413) xor data_in(415) xor data_in(417) xor data_in(423) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(430) xor data_in(431) xor data_in(432) xor data_in(433) xor data_in(435) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(441) xor data_in(443) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(449) xor data_in(450) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(456) xor data_in(460) xor data_in(462) xor data_in(465) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(472) xor data_in(474) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(481) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(496) xor data_in(498) xor data_in(502) xor data_in(503) xor data_in(507) xor data_in(508) xor data_in(509);
    crc_out(49) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(3) xor crc_in(10) xor crc_in(11) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(18) xor crc_in(19) xor crc_in(20) xor crc_in(21) xor crc_in(24) xor crc_in(25) xor crc_in(33) xor crc_in(35) xor crc_in(36) xor crc_in(37) xor crc_in(43) xor crc_in(48) xor crc_in(49) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(59) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(10) xor data_in(11) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(24) xor data_in(25) xor data_in(33) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(43) xor data_in(48) xor data_in(49) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(64) xor data_in(65) xor data_in(67) xor data_in(68) xor data_in(71) xor data_in(72) xor data_in(75) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(90) xor data_in(91) xor data_in(93) xor data_in(98) xor data_in(99) xor data_in(100) xor data_in(103) xor data_in(107) xor data_in(108) xor data_in(109) xor data_in(111) xor data_in(115) xor data_in(117) xor data_in(119) xor data_in(120) xor data_in(126) xor data_in(128) xor data_in(131) xor data_in(132) xor data_in(134) xor data_in(135) xor data_in(138) xor data_in(141) xor data_in(142) xor data_in(143) xor data_in(144) xor data_in(146) xor data_in(149) xor data_in(151) xor data_in(152) xor data_in(154) xor data_in(155) xor data_in(156) xor data_in(158) xor data_in(160) xor data_in(161) xor data_in(162) xor data_in(167) xor data_in(168) xor data_in(170) xor data_in(171) xor data_in(175) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(182) xor data_in(183) xor data_in(186) xor data_in(187) xor data_in(192) xor data_in(193) xor data_in(195) xor data_in(196) xor data_in(197) xor data_in(200) xor data_in(201) xor data_in(202) xor data_in(209) xor data_in(210) xor data_in(215) xor data_in(217) xor data_in(219) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(223) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(238) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(242) xor data_in(243) xor data_in(247) xor data_in(248) xor data_in(250) xor data_in(251) xor data_in(252) xor data_in(254) xor data_in(257) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(268) xor data_in(269) xor data_in(271) xor data_in(272) xor data_in(278) xor data_in(280) xor data_in(282) xor data_in(285) xor data_in(287) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(294) xor data_in(295) xor data_in(298) xor data_in(300) xor data_in(301) xor data_in(303) xor data_in(306) xor data_in(307) xor data_in(308) xor data_in(309) xor data_in(310) xor data_in(315) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(323) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(334) xor data_in(335) xor data_in(336) xor data_in(338) xor data_in(339) xor data_in(340) xor data_in(341) xor data_in(344) xor data_in(345) xor data_in(349) xor data_in(352) xor data_in(355) xor data_in(360) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(370) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(377) xor data_in(378) xor data_in(380) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(385) xor data_in(386) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(393) xor data_in(394) xor data_in(396) xor data_in(401) xor data_in(402) xor data_in(404) xor data_in(405) xor data_in(409) xor data_in(410) xor data_in(412) xor data_in(414) xor data_in(416) xor data_in(418) xor data_in(424) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(429) xor data_in(431) xor data_in(432) xor data_in(433) xor data_in(434) xor data_in(436) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(442) xor data_in(444) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(450) xor data_in(451) xor data_in(454) xor data_in(455) xor data_in(456) xor data_in(457) xor data_in(461) xor data_in(463) xor data_in(466) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(471) xor data_in(473) xor data_in(475) xor data_in(478) xor data_in(479) xor data_in(480) xor data_in(482) xor data_in(488) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(497) xor data_in(499) xor data_in(503) xor data_in(504) xor data_in(508) xor data_in(509) xor data_in(510);
    crc_out(50) <= crc_in(1) xor crc_in(2) xor crc_in(3) xor crc_in(4) xor crc_in(11) xor crc_in(12) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(17) xor crc_in(19) xor crc_in(20) xor crc_in(21) xor crc_in(22) xor crc_in(25) xor crc_in(26) xor crc_in(34) xor crc_in(36) xor crc_in(37) xor crc_in(38) xor crc_in(44) xor crc_in(49) xor crc_in(50) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(56) xor crc_in(57) xor crc_in(60) xor crc_in(61) xor crc_in(62) xor crc_in(63) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(25) xor data_in(26) xor data_in(34) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(44) xor data_in(49) xor data_in(50) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63) xor data_in(64) xor data_in(65) xor data_in(66) xor data_in(68) xor data_in(69) xor data_in(72) xor data_in(73) xor data_in(76) xor data_in(80) xor data_in(81) xor data_in(82) xor data_in(86) xor data_in(87) xor data_in(88) xor data_in(91) xor data_in(92) xor data_in(94) xor data_in(99) xor data_in(100) xor data_in(101) xor data_in(104) xor data_in(108) xor data_in(109) xor data_in(110) xor data_in(112) xor data_in(116) xor data_in(118) xor data_in(120) xor data_in(121) xor data_in(127) xor data_in(129) xor data_in(132) xor data_in(133) xor data_in(135) xor data_in(136) xor data_in(139) xor data_in(142) xor data_in(143) xor data_in(144) xor data_in(145) xor data_in(147) xor data_in(150) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(159) xor data_in(161) xor data_in(162) xor data_in(163) xor data_in(168) xor data_in(169) xor data_in(171) xor data_in(172) xor data_in(176) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(183) xor data_in(184) xor data_in(187) xor data_in(188) xor data_in(193) xor data_in(194) xor data_in(196) xor data_in(197) xor data_in(198) xor data_in(201) xor data_in(202) xor data_in(203) xor data_in(210) xor data_in(211) xor data_in(216) xor data_in(218) xor data_in(220) xor data_in(221) xor data_in(222) xor data_in(223) xor data_in(224) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(242) xor data_in(243) xor data_in(244) xor data_in(248) xor data_in(249) xor data_in(251) xor data_in(252) xor data_in(253) xor data_in(255) xor data_in(258) xor data_in(260) xor data_in(261) xor data_in(262) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(273) xor data_in(279) xor data_in(281) xor data_in(283) xor data_in(286) xor data_in(288) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(295) xor data_in(296) xor data_in(299) xor data_in(301) xor data_in(302) xor data_in(304) xor data_in(307) xor data_in(308) xor data_in(309) xor data_in(310) xor data_in(311) xor data_in(316) xor data_in(318) xor data_in(319) xor data_in(320) xor data_in(321) xor data_in(324) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(335) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(340) xor data_in(341) xor data_in(342) xor data_in(345) xor data_in(346) xor data_in(350) xor data_in(353) xor data_in(356) xor data_in(361) xor data_in(364) xor data_in(365) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(371) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(378) xor data_in(379) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(386) xor data_in(387) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(394) xor data_in(395) xor data_in(397) xor data_in(402) xor data_in(403) xor data_in(405) xor data_in(406) xor data_in(410) xor data_in(411) xor data_in(413) xor data_in(415) xor data_in(417) xor data_in(419) xor data_in(425) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(429) xor data_in(430) xor data_in(432) xor data_in(433) xor data_in(434) xor data_in(435) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(440) xor data_in(443) xor data_in(445) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(449) xor data_in(451) xor data_in(452) xor data_in(455) xor data_in(456) xor data_in(457) xor data_in(458) xor data_in(462) xor data_in(464) xor data_in(467) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(471) xor data_in(472) xor data_in(474) xor data_in(476) xor data_in(479) xor data_in(480) xor data_in(481) xor data_in(483) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(498) xor data_in(500) xor data_in(504) xor data_in(505) xor data_in(509) xor data_in(510) xor data_in(511);
    crc_out(51) <= crc_in(3) xor crc_in(4) xor crc_in(7) xor crc_in(8) xor crc_in(10) xor crc_in(14) xor crc_in(16) xor crc_in(17) xor crc_in(18) xor crc_in(20) xor crc_in(23) xor crc_in(24) xor crc_in(26) xor crc_in(27) xor crc_in(32) xor crc_in(35) xor crc_in(36) xor crc_in(37) xor crc_in(38) xor crc_in(39) xor crc_in(41) xor crc_in(43) xor crc_in(47) xor crc_in(51) xor crc_in(52) xor crc_in(53) xor crc_in(56) xor crc_in(57) xor crc_in(59) xor crc_in(61) xor crc_in(63) xor data_in(3) xor data_in(4) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(32) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(47) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(56) xor data_in(57) xor data_in(59) xor data_in(61) xor data_in(63) xor data_in(64) xor data_in(65) xor data_in(66) xor data_in(67) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(76) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(85) xor data_in(86) xor data_in(88) xor data_in(89) xor data_in(93) xor data_in(100) xor data_in(101) xor data_in(103) xor data_in(104) xor data_in(105) xor data_in(108) xor data_in(109) xor data_in(114) xor data_in(117) xor data_in(120) xor data_in(121) xor data_in(123) xor data_in(124) xor data_in(126) xor data_in(128) xor data_in(129) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(138) xor data_in(139) xor data_in(141) xor data_in(142) xor data_in(144) xor data_in(145) xor data_in(148) xor data_in(150) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(162) xor data_in(163) xor data_in(165) xor data_in(166) xor data_in(167) xor data_in(168) xor data_in(169) xor data_in(171) xor data_in(172) xor data_in(173) xor data_in(175) xor data_in(176) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(185) xor data_in(186) xor data_in(188) xor data_in(189) xor data_in(190) xor data_in(195) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(202) xor data_in(203) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(208) xor data_in(214) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(219) xor data_in(221) xor data_in(222) xor data_in(226) xor data_in(228) xor data_in(229) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(243) xor data_in(244) xor data_in(249) xor data_in(250) xor data_in(253) xor data_in(256) xor data_in(258) xor data_in(259) xor data_in(261) xor data_in(264) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(274) xor data_in(275) xor data_in(276) xor data_in(278) xor data_in(280) xor data_in(281) xor data_in(282) xor data_in(284) xor data_in(288) xor data_in(289) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(295) xor data_in(296) xor data_in(298) xor data_in(299) xor data_in(304) xor data_in(305) xor data_in(308) xor data_in(310) xor data_in(311) xor data_in(312) xor data_in(313) xor data_in(314) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(326) xor data_in(327) xor data_in(330) xor data_in(331) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(341) xor data_in(342) xor data_in(344) xor data_in(345) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(351) xor data_in(352) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(358) xor data_in(363) xor data_in(364) xor data_in(365) xor data_in(366) xor data_in(369) xor data_in(370) xor data_in(373) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(383) xor data_in(384) xor data_in(396) xor data_in(397) xor data_in(400) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(411) xor data_in(413) xor data_in(414) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(421) xor data_in(423) xor data_in(424) xor data_in(426) xor data_in(427) xor data_in(428) xor data_in(433) xor data_in(436) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(444) xor data_in(446) xor data_in(447) xor data_in(448) xor data_in(450) xor data_in(454) xor data_in(456) xor data_in(457) xor data_in(458) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(465) xor data_in(466) xor data_in(468) xor data_in(469) xor data_in(472) xor data_in(473) xor data_in(474) xor data_in(478) xor data_in(480) xor data_in(481) xor data_in(482) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(490) xor data_in(492) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(498) xor data_in(501) xor data_in(503) xor data_in(504) xor data_in(508) xor data_in(511);
    crc_out(52) <= crc_in(2) xor crc_in(4) xor crc_in(7) xor crc_in(9) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(17) xor crc_in(18) xor crc_in(19) xor crc_in(22) xor crc_in(25) xor crc_in(27) xor crc_in(28) xor crc_in(32) xor crc_in(33) xor crc_in(37) xor crc_in(38) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(47) xor crc_in(48) xor crc_in(50) xor crc_in(55) xor crc_in(57) xor crc_in(59) xor crc_in(60) xor data_in(2) xor data_in(4) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(22) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(32) xor data_in(33) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(48) xor data_in(50) xor data_in(55) xor data_in(57) xor data_in(59) xor data_in(60) xor data_in(64) xor data_in(65) xor data_in(66) xor data_in(67) xor data_in(68) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(73) xor data_in(76) xor data_in(78) xor data_in(81) xor data_in(83) xor data_in(85) xor data_in(89) xor data_in(90) xor data_in(92) xor data_in(94) xor data_in(95) xor data_in(101) xor data_in(103) xor data_in(105) xor data_in(106) xor data_in(108) xor data_in(109) xor data_in(111) xor data_in(113) xor data_in(114) xor data_in(115) xor data_in(118) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(123) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(141) xor data_in(145) xor data_in(149) xor data_in(150) xor data_in(152) xor data_in(153) xor data_in(155) xor data_in(157) xor data_in(158) xor data_in(160) xor data_in(163) xor data_in(165) xor data_in(169) xor data_in(171) xor data_in(172) xor data_in(173) xor data_in(174) xor data_in(175) xor data_in(178) xor data_in(180) xor data_in(182) xor data_in(184) xor data_in(187) xor data_in(189) xor data_in(191) xor data_in(194) xor data_in(196) xor data_in(197) xor data_in(199) xor data_in(201) xor data_in(203) xor data_in(205) xor data_in(209) xor data_in(211) xor data_in(212) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(219) xor data_in(220) xor data_in(222) xor data_in(224) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(239) xor data_in(240) xor data_in(241) xor data_in(244) xor data_in(250) xor data_in(251) xor data_in(252) xor data_in(257) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(263) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(277) xor data_in(278) xor data_in(279) xor data_in(282) xor data_in(283) xor data_in(285) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(296) xor data_in(298) xor data_in(302) xor data_in(303) xor data_in(304) xor data_in(305) xor data_in(306) xor data_in(311) xor data_in(312) xor data_in(315) xor data_in(319) xor data_in(322) xor data_in(324) xor data_in(325) xor data_in(326) xor data_in(328) xor data_in(330) xor data_in(333) xor data_in(334) xor data_in(337) xor data_in(339) xor data_in(342) xor data_in(344) xor data_in(350) xor data_in(354) xor data_in(358) xor data_in(359) xor data_in(362) xor data_in(363) xor data_in(365) xor data_in(366) xor data_in(368) xor data_in(370) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(380) xor data_in(382) xor data_in(384) xor data_in(387) xor data_in(388) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(395) xor data_in(400) xor data_in(401) xor data_in(404) xor data_in(406) xor data_in(407) xor data_in(410) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(425) xor data_in(427) xor data_in(428) xor data_in(430) xor data_in(431) xor data_in(435) xor data_in(437) xor data_in(438) xor data_in(439) xor data_in(441) xor data_in(443) xor data_in(445) xor data_in(447) xor data_in(448) xor data_in(451) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(457) xor data_in(458) xor data_in(460) xor data_in(467) xor data_in(469) xor data_in(471) xor data_in(473) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(481) xor data_in(482) xor data_in(483) xor data_in(484) xor data_in(486) xor data_in(489) xor data_in(495) xor data_in(497) xor data_in(498) xor data_in(502) xor data_in(503) xor data_in(506) xor data_in(508) xor data_in(509) xor data_in(510);
    crc_out(53) <= crc_in(0) xor crc_in(3) xor crc_in(5) xor crc_in(8) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(18) xor crc_in(19) xor crc_in(20) xor crc_in(23) xor crc_in(26) xor crc_in(28) xor crc_in(29) xor crc_in(33) xor crc_in(34) xor crc_in(38) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(48) xor crc_in(49) xor crc_in(51) xor crc_in(56) xor crc_in(58) xor crc_in(60) xor crc_in(61) xor data_in(0) xor data_in(3) xor data_in(5) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(23) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(33) xor data_in(34) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(48) xor data_in(49) xor data_in(51) xor data_in(56) xor data_in(58) xor data_in(60) xor data_in(61) xor data_in(65) xor data_in(66) xor data_in(67) xor data_in(68) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(74) xor data_in(77) xor data_in(79) xor data_in(82) xor data_in(84) xor data_in(86) xor data_in(90) xor data_in(91) xor data_in(93) xor data_in(95) xor data_in(96) xor data_in(102) xor data_in(104) xor data_in(106) xor data_in(107) xor data_in(109) xor data_in(110) xor data_in(112) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(119) xor data_in(120) xor data_in(121) xor data_in(122) xor data_in(124) xor data_in(126) xor data_in(127) xor data_in(128) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(142) xor data_in(146) xor data_in(150) xor data_in(151) xor data_in(153) xor data_in(154) xor data_in(156) xor data_in(158) xor data_in(159) xor data_in(161) xor data_in(164) xor data_in(166) xor data_in(170) xor data_in(172) xor data_in(173) xor data_in(174) xor data_in(175) xor data_in(176) xor data_in(179) xor data_in(181) xor data_in(183) xor data_in(185) xor data_in(188) xor data_in(190) xor data_in(192) xor data_in(195) xor data_in(197) xor data_in(198) xor data_in(200) xor data_in(202) xor data_in(204) xor data_in(206) xor data_in(210) xor data_in(212) xor data_in(213) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(218) xor data_in(220) xor data_in(221) xor data_in(223) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(240) xor data_in(241) xor data_in(242) xor data_in(245) xor data_in(251) xor data_in(252) xor data_in(253) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(275) xor data_in(278) xor data_in(279) xor data_in(280) xor data_in(283) xor data_in(284) xor data_in(286) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(295) xor data_in(297) xor data_in(299) xor data_in(303) xor data_in(304) xor data_in(305) xor data_in(306) xor data_in(307) xor data_in(312) xor data_in(313) xor data_in(316) xor data_in(320) xor data_in(323) xor data_in(325) xor data_in(326) xor data_in(327) xor data_in(329) xor data_in(331) xor data_in(334) xor data_in(335) xor data_in(338) xor data_in(340) xor data_in(343) xor data_in(345) xor data_in(351) xor data_in(355) xor data_in(359) xor data_in(360) xor data_in(363) xor data_in(364) xor data_in(366) xor data_in(367) xor data_in(369) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(375) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(380) xor data_in(381) xor data_in(383) xor data_in(385) xor data_in(388) xor data_in(389) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(396) xor data_in(401) xor data_in(402) xor data_in(405) xor data_in(407) xor data_in(408) xor data_in(411) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(418) xor data_in(419) xor data_in(422) xor data_in(423) xor data_in(424) xor data_in(426) xor data_in(428) xor data_in(429) xor data_in(431) xor data_in(432) xor data_in(436) xor data_in(438) xor data_in(439) xor data_in(440) xor data_in(442) xor data_in(444) xor data_in(446) xor data_in(448) xor data_in(449) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(455) xor data_in(456) xor data_in(458) xor data_in(459) xor data_in(461) xor data_in(468) xor data_in(470) xor data_in(472) xor data_in(474) xor data_in(478) xor data_in(479) xor data_in(480) xor data_in(482) xor data_in(483) xor data_in(484) xor data_in(485) xor data_in(487) xor data_in(490) xor data_in(496) xor data_in(498) xor data_in(499) xor data_in(503) xor data_in(504) xor data_in(507) xor data_in(509) xor data_in(510) xor data_in(511);
    crc_out(54) <= crc_in(0) xor crc_in(1) xor crc_in(2) xor crc_in(4) xor crc_in(5) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(10) xor crc_in(11) xor crc_in(16) xor crc_in(19) xor crc_in(20) xor crc_in(22) xor crc_in(27) xor crc_in(29) xor crc_in(30) xor crc_in(32) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(39) xor crc_in(40) xor crc_in(42) xor crc_in(44) xor crc_in(46) xor crc_in(49) xor crc_in(53) xor crc_in(54) xor crc_in(55) xor crc_in(57) xor crc_in(58) xor crc_in(61) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(16) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(39) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(46) xor data_in(49) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(57) xor data_in(58) xor data_in(61) xor data_in(66) xor data_in(67) xor data_in(68) xor data_in(73) xor data_in(74) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(79) xor data_in(82) xor data_in(86) xor data_in(91) xor data_in(94) xor data_in(95) xor data_in(96) xor data_in(97) xor data_in(102) xor data_in(104) xor data_in(105) xor data_in(107) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(119) xor data_in(121) xor data_in(124) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(128) xor data_in(130) xor data_in(132) xor data_in(134) xor data_in(135) xor data_in(141) xor data_in(142) xor data_in(146) xor data_in(147) xor data_in(150) xor data_in(156) xor data_in(158) xor data_in(159) xor data_in(162) xor data_in(164) xor data_in(166) xor data_in(168) xor data_in(170) xor data_in(173) xor data_in(174) xor data_in(178) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(189) xor data_in(190) xor data_in(191) xor data_in(193) xor data_in(194) xor data_in(196) xor data_in(197) xor data_in(198) xor data_in(199) xor data_in(200) xor data_in(201) xor data_in(203) xor data_in(204) xor data_in(206) xor data_in(208) xor data_in(212) xor data_in(213) xor data_in(217) xor data_in(219) xor data_in(221) xor data_in(222) xor data_in(223) xor data_in(225) xor data_in(227) xor data_in(231) xor data_in(232) xor data_in(238) xor data_in(241) xor data_in(243) xor data_in(245) xor data_in(246) xor data_in(253) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(263) xor data_in(264) xor data_in(265) xor data_in(270) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(275) xor data_in(278) xor data_in(279) xor data_in(280) xor data_in(284) xor data_in(285) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(296) xor data_in(297) xor data_in(299) xor data_in(302) xor data_in(303) xor data_in(305) xor data_in(306) xor data_in(307) xor data_in(308) xor data_in(309) xor data_in(317) xor data_in(318) xor data_in(320) xor data_in(321) xor data_in(323) xor data_in(324) xor data_in(325) xor data_in(328) xor data_in(331) xor data_in(333) xor data_in(334) xor data_in(335) xor data_in(336) xor data_in(338) xor data_in(340) xor data_in(341) xor data_in(343) xor data_in(345) xor data_in(348) xor data_in(349) xor data_in(353) xor data_in(355) xor data_in(357) xor data_in(358) xor data_in(360) xor data_in(361) xor data_in(362) xor data_in(363) xor data_in(365) xor data_in(370) xor data_in(374) xor data_in(375) xor data_in(376) xor data_in(378) xor data_in(381) xor data_in(384) xor data_in(385) xor data_in(386) xor data_in(387) xor data_in(388) xor data_in(389) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(394) xor data_in(398) xor data_in(400) xor data_in(402) xor data_in(403) xor data_in(405) xor data_in(406) xor data_in(413) xor data_in(415) xor data_in(418) xor data_in(421) xor data_in(425) xor data_in(427) xor data_in(431) xor data_in(432) xor data_in(433) xor data_in(434) xor data_in(435) xor data_in(437) xor data_in(438) xor data_in(440) xor data_in(441) xor data_in(442) xor data_in(443) xor data_in(445) xor data_in(447) xor data_in(450) xor data_in(452) xor data_in(455) xor data_in(456) xor data_in(457) xor data_in(461) xor data_in(463) xor data_in(466) xor data_in(469) xor data_in(470) xor data_in(473) xor data_in(474) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(480) xor data_in(481) xor data_in(483) xor data_in(485) xor data_in(487) xor data_in(493) xor data_in(496) xor data_in(497) xor data_in(498) xor data_in(500) xor data_in(503) xor data_in(506) xor data_in(511);
    crc_out(55) <= crc_in(0) xor crc_in(1) xor crc_in(3) xor crc_in(6) xor crc_in(9) xor crc_in(11) xor crc_in(13) xor crc_in(14) xor crc_in(15) xor crc_in(17) xor crc_in(20) xor crc_in(22) xor crc_in(23) xor crc_in(24) xor crc_in(28) xor crc_in(30) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(35) xor crc_in(37) xor crc_in(40) xor crc_in(52) xor crc_in(53) xor crc_in(56) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(6) xor data_in(9) xor data_in(11) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(35) xor data_in(37) xor data_in(40) xor data_in(52) xor data_in(53) xor data_in(56) xor data_in(67) xor data_in(68) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(75) xor data_in(79) xor data_in(82) xor data_in(85) xor data_in(86) xor data_in(96) xor data_in(97) xor data_in(98) xor data_in(102) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(110) xor data_in(111) xor data_in(113) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(127) xor data_in(128) xor data_in(130) xor data_in(131) xor data_in(132) xor data_in(133) xor data_in(135) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(146) xor data_in(147) xor data_in(148) xor data_in(150) xor data_in(152) xor data_in(154) xor data_in(155) xor data_in(156) xor data_in(158) xor data_in(159) xor data_in(163) xor data_in(164) xor data_in(166) xor data_in(168) xor data_in(169) xor data_in(170) xor data_in(174) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(180) xor data_in(184) xor data_in(186) xor data_in(191) xor data_in(192) xor data_in(195) xor data_in(198) xor data_in(199) xor data_in(201) xor data_in(202) xor data_in(206) xor data_in(208) xor data_in(209) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(216) xor data_in(220) xor data_in(222) xor data_in(225) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(244) xor data_in(245) xor data_in(246) xor data_in(247) xor data_in(252) xor data_in(258) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(263) xor data_in(265) xor data_in(267) xor data_in(268) xor data_in(269) xor data_in(271) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(278) xor data_in(279) xor data_in(280) xor data_in(285) xor data_in(286) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(293) xor data_in(294) xor data_in(299) xor data_in(302) xor data_in(306) xor data_in(307) xor data_in(308) xor data_in(310) xor data_in(313) xor data_in(314) xor data_in(319) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(324) xor data_in(327) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(333) xor data_in(335) xor data_in(336) xor data_in(337) xor data_in(338) xor data_in(340) xor data_in(341) xor data_in(342) xor data_in(343) xor data_in(345) xor data_in(348) xor data_in(350) xor data_in(352) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(357) xor data_in(359) xor data_in(361) xor data_in(366) xor data_in(367) xor data_in(368) xor data_in(371) xor data_in(372) xor data_in(373) xor data_in(375) xor data_in(376) xor data_in(377) xor data_in(380) xor data_in(386) xor data_in(389) xor data_in(390) xor data_in(397) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(417) xor data_in(420) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(424) xor data_in(426) xor data_in(428) xor data_in(429) xor data_in(430) xor data_in(431) xor data_in(432) xor data_in(433) xor data_in(436) xor data_in(441) xor data_in(443) xor data_in(444) xor data_in(446) xor data_in(448) xor data_in(449) xor data_in(451) xor data_in(452) xor data_in(454) xor data_in(456) xor data_in(457) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(463) xor data_in(464) xor data_in(466) xor data_in(467) xor data_in(477) xor data_in(479) xor data_in(480) xor data_in(481) xor data_in(482) xor data_in(487) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(496) xor data_in(497) xor data_in(501) xor data_in(503) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(510);
    crc_out(56) <= crc_in(1) xor crc_in(2) xor crc_in(4) xor crc_in(7) xor crc_in(10) xor crc_in(12) xor crc_in(14) xor crc_in(15) xor crc_in(16) xor crc_in(18) xor crc_in(21) xor crc_in(23) xor crc_in(24) xor crc_in(25) xor crc_in(29) xor crc_in(31) xor crc_in(32) xor crc_in(33) xor crc_in(34) xor crc_in(36) xor crc_in(38) xor crc_in(41) xor crc_in(53) xor crc_in(54) xor crc_in(57) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(7) xor data_in(10) xor data_in(12) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(36) xor data_in(38) xor data_in(41) xor data_in(53) xor data_in(54) xor data_in(57) xor data_in(68) xor data_in(69) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(76) xor data_in(80) xor data_in(83) xor data_in(86) xor data_in(87) xor data_in(97) xor data_in(98) xor data_in(99) xor data_in(103) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(111) xor data_in(112) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(120) xor data_in(124) xor data_in(125) xor data_in(126) xor data_in(128) xor data_in(129) xor data_in(131) xor data_in(132) xor data_in(133) xor data_in(134) xor data_in(136) xor data_in(138) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(142) xor data_in(147) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(153) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(159) xor data_in(160) xor data_in(164) xor data_in(165) xor data_in(167) xor data_in(169) xor data_in(170) xor data_in(171) xor data_in(175) xor data_in(177) xor data_in(178) xor data_in(179) xor data_in(181) xor data_in(185) xor data_in(187) xor data_in(192) xor data_in(193) xor data_in(196) xor data_in(199) xor data_in(200) xor data_in(202) xor data_in(203) xor data_in(207) xor data_in(209) xor data_in(210) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(217) xor data_in(221) xor data_in(223) xor data_in(226) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(245) xor data_in(246) xor data_in(247) xor data_in(248) xor data_in(253) xor data_in(259) xor data_in(260) xor data_in(261) xor data_in(262) xor data_in(264) xor data_in(266) xor data_in(268) xor data_in(269) xor data_in(270) xor data_in(272) xor data_in(273) xor data_in(274) xor data_in(275) xor data_in(279) xor data_in(280) xor data_in(281) xor data_in(286) xor data_in(287) xor data_in(288) xor data_in(289) xor data_in(290) xor data_in(291) xor data_in(294) xor data_in(295) xor data_in(300) xor data_in(303) xor data_in(307) xor data_in(308) xor data_in(309) xor data_in(311) xor data_in(314) xor data_in(315) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(324) xor data_in(325) xor data_in(328) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(334) xor data_in(336) xor data_in(337) xor data_in(338) xor data_in(339) xor data_in(341) xor data_in(342) xor data_in(343) xor data_in(344) xor data_in(346) xor data_in(349) xor data_in(351) xor data_in(353) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(358) xor data_in(360) xor data_in(362) xor data_in(367) xor data_in(368) xor data_in(369) xor data_in(372) xor data_in(373) xor data_in(374) xor data_in(376) xor data_in(377) xor data_in(378) xor data_in(381) xor data_in(387) xor data_in(390) xor data_in(391) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(402) xor data_in(404) xor data_in(405) xor data_in(406) xor data_in(407) xor data_in(408) xor data_in(409) xor data_in(410) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(418) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(424) xor data_in(425) xor data_in(427) xor data_in(429) xor data_in(430) xor data_in(431) xor data_in(432) xor data_in(433) xor data_in(434) xor data_in(437) xor data_in(442) xor data_in(444) xor data_in(445) xor data_in(447) xor data_in(449) xor data_in(450) xor data_in(452) xor data_in(453) xor data_in(455) xor data_in(457) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(464) xor data_in(465) xor data_in(467) xor data_in(468) xor data_in(478) xor data_in(480) xor data_in(481) xor data_in(482) xor data_in(483) xor data_in(488) xor data_in(492) xor data_in(494) xor data_in(495) xor data_in(497) xor data_in(498) xor data_in(502) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(509) xor data_in(511);
    crc_out(57) <= crc_in(0) xor crc_in(3) xor crc_in(7) xor crc_in(10) xor crc_in(11) xor crc_in(12) xor crc_in(14) xor crc_in(16) xor crc_in(17) xor crc_in(19) xor crc_in(21) xor crc_in(25) xor crc_in(26) xor crc_in(30) xor crc_in(33) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(37) xor crc_in(39) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(45) xor crc_in(47) xor crc_in(50) xor crc_in(52) xor crc_in(53) xor crc_in(59) xor crc_in(62) xor data_in(0) xor data_in(3) xor data_in(7) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(21) xor data_in(25) xor data_in(26) xor data_in(30) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(45) xor data_in(47) xor data_in(50) xor data_in(52) xor data_in(53) xor data_in(59) xor data_in(62) xor data_in(71) xor data_in(73) xor data_in(76) xor data_in(78) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(88) xor data_in(92) xor data_in(95) xor data_in(98) xor data_in(99) xor data_in(100) xor data_in(102) xor data_in(103) xor data_in(106) xor data_in(107) xor data_in(110) xor data_in(111) xor data_in(112) xor data_in(114) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(127) xor data_in(133) xor data_in(134) xor data_in(135) xor data_in(136) xor data_in(138) xor data_in(146) xor data_in(148) xor data_in(149) xor data_in(151) xor data_in(155) xor data_in(161) xor data_in(164) xor data_in(167) xor data_in(172) xor data_in(175) xor data_in(177) xor data_in(180) xor data_in(181) xor data_in(184) xor data_in(188) xor data_in(190) xor data_in(193) xor data_in(201) xor data_in(203) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(210) xor data_in(212) xor data_in(213) xor data_in(215) xor data_in(216) xor data_in(222) xor data_in(223) xor data_in(225) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(234) xor data_in(235) xor data_in(238) xor data_in(242) xor data_in(245) xor data_in(246) xor data_in(247) xor data_in(248) xor data_in(249) xor data_in(252) xor data_in(258) xor data_in(260) xor data_in(261) xor data_in(264) xor data_in(265) xor data_in(266) xor data_in(268) xor data_in(270) xor data_in(271) xor data_in(273) xor data_in(274) xor data_in(278) xor data_in(280) xor data_in(282) xor data_in(289) xor data_in(290) xor data_in(292) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(308) xor data_in(310) xor data_in(312) xor data_in(313) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(318) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(324) xor data_in(327) xor data_in(329) xor data_in(330) xor data_in(334) xor data_in(335) xor data_in(337) xor data_in(342) xor data_in(346) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(353) xor data_in(354) xor data_in(358) xor data_in(359) xor data_in(361) xor data_in(362) xor data_in(364) xor data_in(367) xor data_in(369) xor data_in(370) xor data_in(372) xor data_in(374) xor data_in(375) xor data_in(377) xor data_in(378) xor data_in(380) xor data_in(385) xor data_in(387) xor data_in(393) xor data_in(395) xor data_in(397) xor data_in(398) xor data_in(399) xor data_in(401) xor data_in(402) xor data_in(403) xor data_in(406) xor data_in(407) xor data_in(410) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(417) xor data_in(420) xor data_in(421) xor data_in(422) xor data_in(425) xor data_in(426) xor data_in(428) xor data_in(429) xor data_in(432) xor data_in(433) xor data_in(439) xor data_in(442) xor data_in(443) xor data_in(445) xor data_in(446) xor data_in(448) xor data_in(449) xor data_in(450) xor data_in(451) xor data_in(452) xor data_in(456) xor data_in(458) xor data_in(465) xor data_in(468) xor data_in(469) xor data_in(470) xor data_in(471) xor data_in(474) xor data_in(475) xor data_in(477) xor data_in(478) xor data_in(479) xor data_in(481) xor data_in(482) xor data_in(483) xor data_in(486) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(491) xor data_in(495) xor data_in(504) xor data_in(506) xor data_in(507) xor data_in(509);
    crc_out(58) <= crc_in(1) xor crc_in(4) xor crc_in(8) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(15) xor crc_in(17) xor crc_in(18) xor crc_in(20) xor crc_in(22) xor crc_in(26) xor crc_in(27) xor crc_in(31) xor crc_in(34) xor crc_in(35) xor crc_in(36) xor crc_in(37) xor crc_in(38) xor crc_in(40) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(46) xor crc_in(48) xor crc_in(51) xor crc_in(53) xor crc_in(54) xor crc_in(60) xor crc_in(63) xor data_in(1) xor data_in(4) xor data_in(8) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(22) xor data_in(26) xor data_in(27) xor data_in(31) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(48) xor data_in(51) xor data_in(53) xor data_in(54) xor data_in(60) xor data_in(63) xor data_in(72) xor data_in(74) xor data_in(77) xor data_in(79) xor data_in(80) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(89) xor data_in(93) xor data_in(96) xor data_in(99) xor data_in(100) xor data_in(101) xor data_in(103) xor data_in(104) xor data_in(107) xor data_in(108) xor data_in(111) xor data_in(112) xor data_in(113) xor data_in(115) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(126) xor data_in(128) xor data_in(134) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(139) xor data_in(147) xor data_in(149) xor data_in(150) xor data_in(152) xor data_in(156) xor data_in(162) xor data_in(165) xor data_in(168) xor data_in(173) xor data_in(176) xor data_in(178) xor data_in(181) xor data_in(182) xor data_in(185) xor data_in(189) xor data_in(191) xor data_in(194) xor data_in(202) xor data_in(204) xor data_in(206) xor data_in(207) xor data_in(208) xor data_in(211) xor data_in(213) xor data_in(214) xor data_in(216) xor data_in(217) xor data_in(223) xor data_in(224) xor data_in(226) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(235) xor data_in(236) xor data_in(239) xor data_in(243) xor data_in(246) xor data_in(247) xor data_in(248) xor data_in(249) xor data_in(250) xor data_in(253) xor data_in(259) xor data_in(261) xor data_in(262) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(269) xor data_in(271) xor data_in(272) xor data_in(274) xor data_in(275) xor data_in(279) xor data_in(281) xor data_in(283) xor data_in(290) xor data_in(291) xor data_in(293) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(304) xor data_in(309) xor data_in(311) xor data_in(313) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(319) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(325) xor data_in(328) xor data_in(330) xor data_in(331) xor data_in(335) xor data_in(336) xor data_in(338) xor data_in(343) xor data_in(347) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(354) xor data_in(355) xor data_in(359) xor data_in(360) xor data_in(362) xor data_in(363) xor data_in(365) xor data_in(368) xor data_in(370) xor data_in(371) xor data_in(373) xor data_in(375) xor data_in(376) xor data_in(378) xor data_in(379) xor data_in(381) xor data_in(386) xor data_in(388) xor data_in(394) xor data_in(396) xor data_in(398) xor data_in(399) xor data_in(400) xor data_in(402) xor data_in(403) xor data_in(404) xor data_in(407) xor data_in(408) xor data_in(411) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(418) xor data_in(421) xor data_in(422) xor data_in(423) xor data_in(426) xor data_in(427) xor data_in(429) xor data_in(430) xor data_in(433) xor data_in(434) xor data_in(440) xor data_in(443) xor data_in(444) xor data_in(446) xor data_in(447) xor data_in(449) xor data_in(450) xor data_in(451) xor data_in(452) xor data_in(453) xor data_in(457) xor data_in(459) xor data_in(466) xor data_in(469) xor data_in(470) xor data_in(471) xor data_in(472) xor data_in(475) xor data_in(476) xor data_in(478) xor data_in(479) xor data_in(480) xor data_in(482) xor data_in(483) xor data_in(484) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(490) xor data_in(492) xor data_in(496) xor data_in(505) xor data_in(507) xor data_in(508) xor data_in(510);
    crc_out(59) <= crc_in(0) xor crc_in(2) xor crc_in(5) xor crc_in(9) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(16) xor crc_in(18) xor crc_in(19) xor crc_in(21) xor crc_in(23) xor crc_in(27) xor crc_in(28) xor crc_in(32) xor crc_in(35) xor crc_in(36) xor crc_in(37) xor crc_in(38) xor crc_in(39) xor crc_in(41) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(47) xor crc_in(49) xor crc_in(52) xor crc_in(54) xor crc_in(55) xor crc_in(61) xor data_in(0) xor data_in(2) xor data_in(5) xor data_in(9) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(23) xor data_in(27) xor data_in(28) xor data_in(32) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(49) xor data_in(52) xor data_in(54) xor data_in(55) xor data_in(61) xor data_in(64) xor data_in(73) xor data_in(75) xor data_in(78) xor data_in(80) xor data_in(81) xor data_in(82) xor data_in(83) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(87) xor data_in(88) xor data_in(90) xor data_in(94) xor data_in(97) xor data_in(100) xor data_in(101) xor data_in(102) xor data_in(104) xor data_in(105) xor data_in(108) xor data_in(109) xor data_in(112) xor data_in(113) xor data_in(114) xor data_in(116) xor data_in(117) xor data_in(118) xor data_in(119) xor data_in(120) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(126) xor data_in(127) xor data_in(129) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(140) xor data_in(148) xor data_in(150) xor data_in(151) xor data_in(153) xor data_in(157) xor data_in(163) xor data_in(166) xor data_in(169) xor data_in(174) xor data_in(177) xor data_in(179) xor data_in(182) xor data_in(183) xor data_in(186) xor data_in(190) xor data_in(192) xor data_in(195) xor data_in(203) xor data_in(205) xor data_in(207) xor data_in(208) xor data_in(209) xor data_in(212) xor data_in(214) xor data_in(215) xor data_in(217) xor data_in(218) xor data_in(224) xor data_in(225) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(236) xor data_in(237) xor data_in(240) xor data_in(244) xor data_in(247) xor data_in(248) xor data_in(249) xor data_in(250) xor data_in(251) xor data_in(254) xor data_in(260) xor data_in(262) xor data_in(263) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(270) xor data_in(272) xor data_in(273) xor data_in(275) xor data_in(276) xor data_in(280) xor data_in(282) xor data_in(284) xor data_in(291) xor data_in(292) xor data_in(294) xor data_in(298) xor data_in(299) xor data_in(300) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(304) xor data_in(305) xor data_in(310) xor data_in(312) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(320) xor data_in(322) xor data_in(323) xor data_in(324) xor data_in(326) xor data_in(329) xor data_in(331) xor data_in(332) xor data_in(336) xor data_in(337) xor data_in(339) xor data_in(344) xor data_in(348) xor data_in(349) xor data_in(350) xor data_in(351) xor data_in(352) xor data_in(355) xor data_in(356) xor data_in(360) xor data_in(361) xor data_in(363) xor data_in(364) xor data_in(366) xor data_in(369) xor data_in(371) xor data_in(372) xor data_in(374) xor data_in(376) xor data_in(377) xor data_in(379) xor data_in(380) xor data_in(382) xor data_in(387) xor data_in(389) xor data_in(395) xor data_in(397) xor data_in(399) xor data_in(400) xor data_in(401) xor data_in(403) xor data_in(404) xor data_in(405) xor data_in(408) xor data_in(409) xor data_in(412) xor data_in(413) xor data_in(414) xor data_in(415) xor data_in(416) xor data_in(417) xor data_in(419) xor data_in(422) xor data_in(423) xor data_in(424) xor data_in(427) xor data_in(428) xor data_in(430) xor data_in(431) xor data_in(434) xor data_in(435) xor data_in(441) xor data_in(444) xor data_in(445) xor data_in(447) xor data_in(448) xor data_in(450) xor data_in(451) xor data_in(452) xor data_in(453) xor data_in(454) xor data_in(458) xor data_in(460) xor data_in(467) xor data_in(470) xor data_in(471) xor data_in(472) xor data_in(473) xor data_in(476) xor data_in(477) xor data_in(479) xor data_in(480) xor data_in(481) xor data_in(483) xor data_in(484) xor data_in(485) xor data_in(488) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(493) xor data_in(497) xor data_in(506) xor data_in(508) xor data_in(509) xor data_in(511);
    crc_out(60) <= crc_in(1) xor crc_in(2) xor crc_in(3) xor crc_in(5) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(12) xor crc_in(17) xor crc_in(19) xor crc_in(20) xor crc_in(21) xor crc_in(28) xor crc_in(29) xor crc_in(32) xor crc_in(33) xor crc_in(37) xor crc_in(38) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(46) xor crc_in(47) xor crc_in(48) xor crc_in(52) xor crc_in(54) xor crc_in(56) xor crc_in(58) xor crc_in(59) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(12) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(28) xor data_in(29) xor data_in(32) xor data_in(33) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(52) xor data_in(54) xor data_in(56) xor data_in(58) xor data_in(59) xor data_in(65) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(77) xor data_in(78) xor data_in(80) xor data_in(81) xor data_in(84) xor data_in(88) xor data_in(89) xor data_in(91) xor data_in(92) xor data_in(98) xor data_in(101) xor data_in(104) xor data_in(105) xor data_in(106) xor data_in(108) xor data_in(109) xor data_in(111) xor data_in(115) xor data_in(117) xor data_in(118) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(125) xor data_in(127) xor data_in(128) xor data_in(129) xor data_in(132) xor data_in(140) xor data_in(142) xor data_in(143) xor data_in(146) xor data_in(149) xor data_in(150) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(160) xor data_in(165) xor data_in(166) xor data_in(168) xor data_in(171) xor data_in(176) xor data_in(177) xor data_in(179) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(183) xor data_in(186) xor data_in(187) xor data_in(190) xor data_in(191) xor data_in(193) xor data_in(194) xor data_in(196) xor data_in(197) xor data_in(200) xor data_in(205) xor data_in(207) xor data_in(209) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(219) xor data_in(223) xor data_in(224) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(238) xor data_in(239) xor data_in(241) xor data_in(242) xor data_in(248) xor data_in(249) xor data_in(250) xor data_in(251) xor data_in(254) xor data_in(255) xor data_in(258) xor data_in(261) xor data_in(262) xor data_in(266) xor data_in(271) xor data_in(273) xor data_in(274) xor data_in(275) xor data_in(277) xor data_in(278) xor data_in(283) xor data_in(285) xor data_in(287) xor data_in(288) xor data_in(291) xor data_in(292) xor data_in(293) xor data_in(297) xor data_in(298) xor data_in(301) xor data_in(305) xor data_in(306) xor data_in(309) xor data_in(311) xor data_in(314) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(319) xor data_in(320) xor data_in(321) xor data_in(324) xor data_in(326) xor data_in(331) xor data_in(334) xor data_in(337) xor data_in(339) xor data_in(343) xor data_in(344) xor data_in(346) xor data_in(348) xor data_in(350) xor data_in(351) xor data_in(355) xor data_in(358) xor data_in(361) xor data_in(363) xor data_in(365) xor data_in(368) xor data_in(370) xor data_in(375) xor data_in(377) xor data_in(378) xor data_in(379) xor data_in(381) xor data_in(382) xor data_in(383) xor data_in(385) xor data_in(387) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(395) xor data_in(396) xor data_in(397) xor data_in(401) xor data_in(402) xor data_in(404) xor data_in(406) xor data_in(408) xor data_in(410) xor data_in(412) xor data_in(414) xor data_in(415) xor data_in(418) xor data_in(419) xor data_in(421) xor data_in(425) xor data_in(428) xor data_in(430) xor data_in(432) xor data_in(434) xor data_in(436) xor data_in(438) xor data_in(439) xor data_in(445) xor data_in(446) xor data_in(448) xor data_in(451) xor data_in(455) xor data_in(460) xor data_in(462) xor data_in(463) xor data_in(466) xor data_in(468) xor data_in(470) xor data_in(472) xor data_in(473) xor data_in(475) xor data_in(480) xor data_in(481) xor data_in(482) xor data_in(485) xor data_in(487) xor data_in(488) xor data_in(489) xor data_in(490) xor data_in(492) xor data_in(493) xor data_in(494) xor data_in(496) xor data_in(499) xor data_in(503) xor data_in(504) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(509);
    crc_out(61) <= crc_in(0) xor crc_in(2) xor crc_in(3) xor crc_in(4) xor crc_in(6) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(13) xor crc_in(18) xor crc_in(20) xor crc_in(21) xor crc_in(22) xor crc_in(29) xor crc_in(30) xor crc_in(33) xor crc_in(34) xor crc_in(38) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(47) xor crc_in(48) xor crc_in(49) xor crc_in(53) xor crc_in(55) xor crc_in(57) xor crc_in(59) xor crc_in(60) xor data_in(0) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(13) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(29) xor data_in(30) xor data_in(33) xor data_in(34) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(48) xor data_in(49) xor data_in(53) xor data_in(55) xor data_in(57) xor data_in(59) xor data_in(60) xor data_in(66) xor data_in(70) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(78) xor data_in(79) xor data_in(81) xor data_in(82) xor data_in(85) xor data_in(89) xor data_in(90) xor data_in(92) xor data_in(93) xor data_in(99) xor data_in(102) xor data_in(105) xor data_in(106) xor data_in(107) xor data_in(109) xor data_in(110) xor data_in(112) xor data_in(116) xor data_in(118) xor data_in(119) xor data_in(122) xor data_in(123) xor data_in(124) xor data_in(126) xor data_in(128) xor data_in(129) xor data_in(130) xor data_in(133) xor data_in(141) xor data_in(143) xor data_in(144) xor data_in(147) xor data_in(150) xor data_in(151) xor data_in(156) xor data_in(157) xor data_in(158) xor data_in(161) xor data_in(166) xor data_in(167) xor data_in(169) xor data_in(172) xor data_in(177) xor data_in(178) xor data_in(180) xor data_in(181) xor data_in(182) xor data_in(183) xor data_in(184) xor data_in(187) xor data_in(188) xor data_in(191) xor data_in(192) xor data_in(194) xor data_in(195) xor data_in(197) xor data_in(198) xor data_in(201) xor data_in(206) xor data_in(208) xor data_in(210) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(220) xor data_in(224) xor data_in(225) xor data_in(235) xor data_in(236) xor data_in(237) xor data_in(239) xor data_in(240) xor data_in(242) xor data_in(243) xor data_in(249) xor data_in(250) xor data_in(251) xor data_in(252) xor data_in(255) xor data_in(256) xor data_in(259) xor data_in(262) xor data_in(263) xor data_in(267) xor data_in(272) xor data_in(274) xor data_in(275) xor data_in(276) xor data_in(278) xor data_in(279) xor data_in(284) xor data_in(286) xor data_in(288) xor data_in(289) xor data_in(292) xor data_in(293) xor data_in(294) xor data_in(298) xor data_in(299) xor data_in(302) xor data_in(306) xor data_in(307) xor data_in(310) xor data_in(312) xor data_in(315) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(320) xor data_in(321) xor data_in(322) xor data_in(325) xor data_in(327) xor data_in(332) xor data_in(335) xor data_in(338) xor data_in(340) xor data_in(344) xor data_in(345) xor data_in(347) xor data_in(349) xor data_in(351) xor data_in(352) xor data_in(356) xor data_in(359) xor data_in(362) xor data_in(364) xor data_in(366) xor data_in(369) xor data_in(371) xor data_in(376) xor data_in(378) xor data_in(379) xor data_in(380) xor data_in(382) xor data_in(383) xor data_in(384) xor data_in(386) xor data_in(388) xor data_in(391) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(396) xor data_in(397) xor data_in(398) xor data_in(402) xor data_in(403) xor data_in(405) xor data_in(407) xor data_in(409) xor data_in(411) xor data_in(413) xor data_in(415) xor data_in(416) xor data_in(419) xor data_in(420) xor data_in(422) xor data_in(426) xor data_in(429) xor data_in(431) xor data_in(433) xor data_in(435) xor data_in(437) xor data_in(439) xor data_in(440) xor data_in(446) xor data_in(447) xor data_in(449) xor data_in(452) xor data_in(456) xor data_in(461) xor data_in(463) xor data_in(464) xor data_in(467) xor data_in(469) xor data_in(471) xor data_in(473) xor data_in(474) xor data_in(476) xor data_in(481) xor data_in(482) xor data_in(483) xor data_in(486) xor data_in(488) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(493) xor data_in(494) xor data_in(495) xor data_in(497) xor data_in(500) xor data_in(504) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(509) xor data_in(510);
    crc_out(62) <= crc_in(0) xor crc_in(1) xor crc_in(3) xor crc_in(4) xor crc_in(5) xor crc_in(7) xor crc_in(8) xor crc_in(9) xor crc_in(10) xor crc_in(14) xor crc_in(19) xor crc_in(21) xor crc_in(22) xor crc_in(23) xor crc_in(30) xor crc_in(31) xor crc_in(34) xor crc_in(35) xor crc_in(39) xor crc_in(40) xor crc_in(41) xor crc_in(42) xor crc_in(43) xor crc_in(44) xor crc_in(45) xor crc_in(46) xor crc_in(48) xor crc_in(49) xor crc_in(50) xor crc_in(54) xor crc_in(56) xor crc_in(58) xor crc_in(60) xor crc_in(61) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(14) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(30) xor data_in(31) xor data_in(34) xor data_in(35) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(54) xor data_in(56) xor data_in(58) xor data_in(60) xor data_in(61) xor data_in(67) xor data_in(71) xor data_in(72) xor data_in(73) xor data_in(74) xor data_in(79) xor data_in(80) xor data_in(82) xor data_in(83) xor data_in(86) xor data_in(90) xor data_in(91) xor data_in(93) xor data_in(94) xor data_in(100) xor data_in(103) xor data_in(106) xor data_in(107) xor data_in(108) xor data_in(110) xor data_in(111) xor data_in(113) xor data_in(117) xor data_in(119) xor data_in(120) xor data_in(123) xor data_in(124) xor data_in(125) xor data_in(127) xor data_in(129) xor data_in(130) xor data_in(131) xor data_in(134) xor data_in(142) xor data_in(144) xor data_in(145) xor data_in(148) xor data_in(151) xor data_in(152) xor data_in(157) xor data_in(158) xor data_in(159) xor data_in(162) xor data_in(167) xor data_in(168) xor data_in(170) xor data_in(173) xor data_in(178) xor data_in(179) xor data_in(181) xor data_in(182) xor data_in(183) xor data_in(184) xor data_in(185) xor data_in(188) xor data_in(189) xor data_in(192) xor data_in(193) xor data_in(195) xor data_in(196) xor data_in(198) xor data_in(199) xor data_in(202) xor data_in(207) xor data_in(209) xor data_in(211) xor data_in(212) xor data_in(213) xor data_in(214) xor data_in(215) xor data_in(216) xor data_in(217) xor data_in(221) xor data_in(225) xor data_in(226) xor data_in(236) xor data_in(237) xor data_in(238) xor data_in(240) xor data_in(241) xor data_in(243) xor data_in(244) xor data_in(250) xor data_in(251) xor data_in(252) xor data_in(253) xor data_in(256) xor data_in(257) xor data_in(260) xor data_in(263) xor data_in(264) xor data_in(268) xor data_in(273) xor data_in(275) xor data_in(276) xor data_in(277) xor data_in(279) xor data_in(280) xor data_in(285) xor data_in(287) xor data_in(289) xor data_in(290) xor data_in(293) xor data_in(294) xor data_in(295) xor data_in(299) xor data_in(300) xor data_in(303) xor data_in(307) xor data_in(308) xor data_in(311) xor data_in(313) xor data_in(316) xor data_in(317) xor data_in(318) xor data_in(319) xor data_in(321) xor data_in(322) xor data_in(323) xor data_in(326) xor data_in(328) xor data_in(333) xor data_in(336) xor data_in(339) xor data_in(341) xor data_in(345) xor data_in(346) xor data_in(348) xor data_in(350) xor data_in(352) xor data_in(353) xor data_in(357) xor data_in(360) xor data_in(363) xor data_in(365) xor data_in(367) xor data_in(370) xor data_in(372) xor data_in(377) xor data_in(379) xor data_in(380) xor data_in(381) xor data_in(383) xor data_in(384) xor data_in(385) xor data_in(387) xor data_in(389) xor data_in(392) xor data_in(393) xor data_in(394) xor data_in(395) xor data_in(397) xor data_in(398) xor data_in(399) xor data_in(403) xor data_in(404) xor data_in(406) xor data_in(408) xor data_in(410) xor data_in(412) xor data_in(414) xor data_in(416) xor data_in(417) xor data_in(420) xor data_in(421) xor data_in(423) xor data_in(427) xor data_in(430) xor data_in(432) xor data_in(434) xor data_in(436) xor data_in(438) xor data_in(440) xor data_in(441) xor data_in(447) xor data_in(448) xor data_in(450) xor data_in(453) xor data_in(457) xor data_in(462) xor data_in(464) xor data_in(465) xor data_in(468) xor data_in(470) xor data_in(472) xor data_in(474) xor data_in(475) xor data_in(477) xor data_in(482) xor data_in(483) xor data_in(484) xor data_in(487) xor data_in(489) xor data_in(490) xor data_in(491) xor data_in(492) xor data_in(494) xor data_in(495) xor data_in(496) xor data_in(498) xor data_in(501) xor data_in(505) xor data_in(506) xor data_in(507) xor data_in(508) xor data_in(509) xor data_in(510) xor data_in(511);
    crc_out(63) <= crc_in(1) xor crc_in(4) xor crc_in(6) xor crc_in(7) xor crc_in(9) xor crc_in(11) xor crc_in(12) xor crc_in(13) xor crc_in(14) xor crc_in(20) xor crc_in(21) xor crc_in(23) xor crc_in(31) xor crc_in(35) xor crc_in(40) xor crc_in(42) xor crc_in(44) xor crc_in(46) xor crc_in(49) xor crc_in(51) xor crc_in(52) xor crc_in(53) xor crc_in(54) xor crc_in(57) xor crc_in(58) xor crc_in(61) xor data_in(1) xor data_in(4) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(31) xor data_in(35) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(46) xor data_in(49) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(57) xor data_in(58) xor data_in(61) xor data_in(68) xor data_in(69) xor data_in(70) xor data_in(71) xor data_in(73) xor data_in(75) xor data_in(76) xor data_in(77) xor data_in(78) xor data_in(79) xor data_in(81) xor data_in(82) xor data_in(84) xor data_in(85) xor data_in(86) xor data_in(91) xor data_in(94) xor data_in(101) xor data_in(102) xor data_in(103) xor data_in(107) xor data_in(109) xor data_in(110) xor data_in(112) xor data_in(113) xor data_in(118) xor data_in(119) xor data_in(121) xor data_in(122) xor data_in(123) xor data_in(125) xor data_in(128) xor data_in(129) xor data_in(131) xor data_in(135) xor data_in(136) xor data_in(137) xor data_in(138) xor data_in(139) xor data_in(140) xor data_in(141) xor data_in(142) xor data_in(145) xor data_in(149) xor data_in(150) xor data_in(151) xor data_in(153) xor data_in(154) xor data_in(155) xor data_in(156) xor data_in(157) xor data_in(159) xor data_in(163) xor data_in(164) xor data_in(165) xor data_in(166) xor data_in(167) xor data_in(169) xor data_in(170) xor data_in(174) xor data_in(175) xor data_in(176) xor data_in(177) xor data_in(178) xor data_in(180) xor data_in(181) xor data_in(183) xor data_in(185) xor data_in(189) xor data_in(193) xor data_in(196) xor data_in(199) xor data_in(203) xor data_in(204) xor data_in(205) xor data_in(206) xor data_in(207) xor data_in(210) xor data_in(211) xor data_in(213) xor data_in(215) xor data_in(217) xor data_in(222) xor data_in(223) xor data_in(224) xor data_in(225) xor data_in(227) xor data_in(228) xor data_in(229) xor data_in(230) xor data_in(231) xor data_in(232) xor data_in(233) xor data_in(234) xor data_in(235) xor data_in(236) xor data_in(238) xor data_in(241) xor data_in(244) xor data_in(251) xor data_in(253) xor data_in(257) xor data_in(261) xor data_in(262) xor data_in(263) xor data_in(265) xor data_in(266) xor data_in(267) xor data_in(268) xor data_in(274) xor data_in(275) xor data_in(277) xor data_in(280) xor data_in(286) xor data_in(287) xor data_in(290) xor data_in(294) xor data_in(296) xor data_in(297) xor data_in(298) xor data_in(299) xor data_in(301) xor data_in(302) xor data_in(303) xor data_in(308) xor data_in(312) xor data_in(313) xor data_in(317) xor data_in(319) xor data_in(322) xor data_in(324) xor data_in(325) xor data_in(326) xor data_in(329) xor data_in(330) xor data_in(331) xor data_in(332) xor data_in(333) xor data_in(337) xor data_in(338) xor data_in(339) xor data_in(342) xor data_in(343) xor data_in(344) xor data_in(345) xor data_in(347) xor data_in(348) xor data_in(351) xor data_in(352) xor data_in(354) xor data_in(355) xor data_in(356) xor data_in(357) xor data_in(361) xor data_in(362) xor data_in(363) xor data_in(366) xor data_in(367) xor data_in(371) xor data_in(372) xor data_in(378) xor data_in(379) xor data_in(381) xor data_in(384) xor data_in(386) xor data_in(387) xor data_in(390) xor data_in(391) xor data_in(392) xor data_in(394) xor data_in(396) xor data_in(397) xor data_in(399) xor data_in(404) xor data_in(407) xor data_in(408) xor data_in(411) xor data_in(412) xor data_in(415) xor data_in(416) xor data_in(418) xor data_in(419) xor data_in(420) xor data_in(422) xor data_in(423) xor data_in(428) xor data_in(429) xor data_in(430) xor data_in(433) xor data_in(434) xor data_in(437) xor data_in(438) xor data_in(441) xor data_in(448) xor data_in(451) xor data_in(452) xor data_in(453) xor data_in(458) xor data_in(459) xor data_in(460) xor data_in(461) xor data_in(462) xor data_in(465) xor data_in(469) xor data_in(470) xor data_in(473) xor data_in(474) xor data_in(476) xor data_in(477) xor data_in(483) xor data_in(485) xor data_in(486) xor data_in(487) xor data_in(490) xor data_in(492) xor data_in(495) xor data_in(497) xor data_in(498) xor data_in(502) xor data_in(503) xor data_in(504) xor data_in(505) xor data_in(507) xor data_in(509) xor data_in(511);
end architecture Behavioral;

-------------------------------------------------------------------------------
-- Copyright (C) 2009 OutputLogic.com
-- This source file may be used and distributed without restriction
-- provided that this copyright statement is not removed from the file
-- and that any derivative work contains the original copyright notice
-- and the associated disclaimer.
--
-- THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
-- WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
-------------------------------------------------------------------------------
-- CRC module for data(63:0)
--   lfsr(63:0)=1+x^1+x^4+x^7+x^9+x^10+x^12+x^13+x^17+x^19+x^21+x^22+x^23+x^24+x^27+x^29+x^31+x^32+x^33+x^35+x^37+x^38+x^39+x^40+x^45+x^46+x^47+x^52+x^53+x^54+x^55+x^57+x^62+x^64;
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity crc is
  port ( data_in : in std_logic_vector (63 downto 0);
    crc_en , rst, clk : in std_logic;
    crc_out : out std_logic_vector (63 downto 0));
end crc;

architecture Behavioral of crc is
  signal lfsr_q: std_logic_vector (63 downto 0);
  signal lfsr_c: std_logic_vector (63 downto 0);
begin
    crc_out <= lfsr_q;

    lfsr_c(0) <= lfsr_q(0) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(26) xor lfsr_q(28) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(46) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(63) xor data_in(0) xor data_in(2) xor data_in(4) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(19) xor data_in(21) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(34) xor data_in(35) xor data_in(37) xor data_in(38) xor data_in(41) xor data_in(42) xor data_in(46) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(63);
    lfsr_c(1) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(10) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(24) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(34) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(49) xor lfsr_q(54) xor lfsr_q(58) xor lfsr_q(61) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(10) xor data_in(13) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(24) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(34) xor data_in(36) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(46) xor data_in(47) xor data_in(49) xor data_in(54) xor data_in(58) xor data_in(61) xor data_in(63);
    lfsr_c(2) <= lfsr_q(1) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(11) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(25) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(44) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(50) xor lfsr_q(55) xor lfsr_q(59) xor lfsr_q(62) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(11) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(25) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(35) xor data_in(37) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(47) xor data_in(48) xor data_in(50) xor data_in(55) xor data_in(59) xor data_in(62);
    lfsr_c(3) <= lfsr_q(2) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(12) xor lfsr_q(15) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(26) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(36) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(45) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(51) xor lfsr_q(56) xor lfsr_q(60) xor lfsr_q(63) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(12) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(36) xor data_in(38) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(45) xor data_in(48) xor data_in(49) xor data_in(51) xor data_in(56) xor data_in(60) xor data_in(63);
    lfsr_c(4) <= lfsr_q(0) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(5) xor lfsr_q(14) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(26) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(44) xor lfsr_q(51) xor lfsr_q(53) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(61) xor lfsr_q(63) xor data_in(0) xor data_in(2) xor data_in(3) xor data_in(5) xor data_in(14) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(44) xor data_in(51) xor data_in(53) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(63);
    lfsr_c(5) <= lfsr_q(1) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(6) xor lfsr_q(15) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(45) xor lfsr_q(52) xor lfsr_q(54) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(61) xor lfsr_q(62) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(6) xor data_in(15) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(35) xor data_in(36) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(45) xor data_in(52) xor data_in(54) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62);
    lfsr_c(6) <= lfsr_q(2) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(16) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(46) xor lfsr_q(53) xor lfsr_q(55) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(61) xor lfsr_q(62) xor lfsr_q(63) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(16) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(36) xor data_in(37) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(46) xor data_in(53) xor data_in(55) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(62) xor data_in(63);
    lfsr_c(7) <= lfsr_q(0) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(23) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(33) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(61) xor lfsr_q(62) xor data_in(0) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(9) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(23) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(33) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(47) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(56) xor data_in(58) xor data_in(59) xor data_in(61) xor data_in(62);
    lfsr_c(8) <= lfsr_q(1) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(24) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(34) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(57) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(62) xor lfsr_q(63) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(8) xor data_in(10) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(24) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(34) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(48) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(57) xor data_in(59) xor data_in(60) xor data_in(62) xor data_in(63);
    lfsr_c(9) <= lfsr_q(0) xor lfsr_q(5) xor lfsr_q(8) xor lfsr_q(11) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(18) xor lfsr_q(24) xor lfsr_q(26) xor lfsr_q(28) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(45) xor lfsr_q(48) xor lfsr_q(50) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(59) xor lfsr_q(61) xor data_in(0) xor data_in(5) xor data_in(8) xor data_in(11) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(18) xor data_in(24) xor data_in(26) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(37) xor data_in(38) xor data_in(41) xor data_in(42) xor data_in(45) xor data_in(48) xor data_in(50) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(59) xor data_in(61);
    lfsr_c(10) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(21) xor lfsr_q(24) xor lfsr_q(26) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(37) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(50) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(62) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(7) xor data_in(8) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(21) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(50) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(62) xor data_in(63);
    lfsr_c(11) <= lfsr_q(1) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(5) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(22) xor lfsr_q(25) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(38) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(44) xor lfsr_q(51) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(63) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(5) xor data_in(8) xor data_in(9) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(22) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(51) xor data_in(53) xor data_in(54) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(63);
    lfsr_c(12) <= lfsr_q(0) xor lfsr_q(3) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(33) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(57) xor lfsr_q(61) xor lfsr_q(63) xor data_in(0) xor data_in(3) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(13) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(33) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(42) xor data_in(43) xor data_in(45) xor data_in(46) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(57) xor data_in(61) xor data_in(63);
    lfsr_c(13) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(2) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(11) xor lfsr_q(13) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(28) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(47) xor lfsr_q(49) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(62) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(6) xor data_in(7) xor data_in(11) xor data_in(13) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(35) xor data_in(37) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(47) xor data_in(49) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(59) xor data_in(60) xor data_in(62) xor data_in(63);
    lfsr_c(14) <= lfsr_q(1) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(12) xor lfsr_q(14) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(29) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(36) xor lfsr_q(38) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(48) xor lfsr_q(50) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(60) xor lfsr_q(61) xor lfsr_q(63) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(7) xor data_in(8) xor data_in(12) xor data_in(14) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(36) xor data_in(38) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(48) xor data_in(50) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(60) xor data_in(61) xor data_in(63);
    lfsr_c(15) <= lfsr_q(2) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(30) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(37) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(49) xor lfsr_q(51) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(61) xor lfsr_q(62) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(8) xor data_in(9) xor data_in(13) xor data_in(15) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(30) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(49) xor data_in(51) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(61) xor data_in(62);
    lfsr_c(16) <= lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(31) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(38) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(50) xor lfsr_q(52) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(62) xor lfsr_q(63) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(9) xor data_in(10) xor data_in(14) xor data_in(16) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(31) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(50) xor data_in(52) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(62) xor data_in(63);
    lfsr_c(17) <= lfsr_q(0) xor lfsr_q(2) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(28) xor lfsr_q(32) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(52) xor lfsr_q(57) xor data_in(0) xor data_in(2) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(22) xor data_in(23) xor data_in(28) xor data_in(32) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(52) xor data_in(57);
    lfsr_c(18) <= lfsr_q(1) xor lfsr_q(3) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(29) xor lfsr_q(33) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(53) xor lfsr_q(58) xor data_in(1) xor data_in(3) xor data_in(6) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(23) xor data_in(24) xor data_in(29) xor data_in(33) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(53) xor data_in(58);
    lfsr_c(19) <= lfsr_q(0) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(26) xor lfsr_q(28) xor lfsr_q(30) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(47) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(58) xor lfsr_q(60) xor lfsr_q(63) xor data_in(0) xor data_in(6) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(26) xor data_in(28) xor data_in(30) xor data_in(35) xor data_in(37) xor data_in(39) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(53) xor data_in(54) xor data_in(58) xor data_in(60) xor data_in(63);
    lfsr_c(20) <= lfsr_q(1) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(27) xor lfsr_q(29) xor lfsr_q(31) xor lfsr_q(36) xor lfsr_q(38) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(48) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(59) xor lfsr_q(61) xor data_in(1) xor data_in(7) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(27) xor data_in(29) xor data_in(31) xor data_in(36) xor data_in(38) xor data_in(40) xor data_in(41) xor data_in(43) xor data_in(45) xor data_in(46) xor data_in(48) xor data_in(54) xor data_in(55) xor data_in(59) xor data_in(61);
    lfsr_c(21) <= lfsr_q(0) xor lfsr_q(4) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(12) xor lfsr_q(17) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(26) xor lfsr_q(30) xor lfsr_q(32) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(44) xor lfsr_q(47) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(62) xor lfsr_q(63) xor data_in(0) xor data_in(4) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(17) xor data_in(20) xor data_in(21) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(30) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(38) xor data_in(39) xor data_in(44) xor data_in(47) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(56) xor data_in(58) xor data_in(59) xor data_in(62) xor data_in(63);
    lfsr_c(22) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(22) xor lfsr_q(24) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(31) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(54) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(14) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(22) xor data_in(24) xor data_in(27) xor data_in(28) xor data_in(31) xor data_in(33) xor data_in(34) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(45) xor data_in(46) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(54) xor data_in(56) xor data_in(57) xor data_in(58);
    lfsr_c(23) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(26) xor lfsr_q(29) xor lfsr_q(32) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(43) xor lfsr_q(47) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(55) xor lfsr_q(57) xor lfsr_q(60) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(29) xor data_in(32) xor data_in(39) xor data_in(40) xor data_in(43) xor data_in(47) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(57) xor data_in(60) xor data_in(63);
    lfsr_c(24) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(15) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(22) xor lfsr_q(26) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(30) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(44) xor lfsr_q(46) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(54) xor lfsr_q(56) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(61) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(22) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(37) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(46) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(54) xor data_in(56) xor data_in(59) xor data_in(60) xor data_in(61) xor data_in(63);
    lfsr_c(25) <= lfsr_q(1) xor lfsr_q(2) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(16) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(23) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(31) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(45) xor lfsr_q(47) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(55) xor lfsr_q(57) xor lfsr_q(60) xor lfsr_q(61) xor lfsr_q(62) xor data_in(1) xor data_in(2) xor data_in(6) xor data_in(8) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(23) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(38) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(45) xor data_in(47) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(57) xor data_in(60) xor data_in(61) xor data_in(62);
    lfsr_c(26) <= lfsr_q(2) xor lfsr_q(3) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(24) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(32) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(44) xor lfsr_q(46) xor lfsr_q(48) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(61) xor lfsr_q(62) xor lfsr_q(63) xor data_in(2) xor data_in(3) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(24) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(39) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(46) xor data_in(48) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(56) xor data_in(58) xor data_in(61) xor data_in(62) xor data_in(63);
    lfsr_c(27) <= lfsr_q(0) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(24) xor lfsr_q(26) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(50) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(60) xor lfsr_q(62) xor data_in(0) xor data_in(2) xor data_in(3) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(24) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(40) xor data_in(42) xor data_in(43) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(50) xor data_in(54) xor data_in(55) xor data_in(57) xor data_in(58) xor data_in(60) xor data_in(62);
    lfsr_c(28) <= lfsr_q(1) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(25) xor lfsr_q(27) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(51) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(61) xor lfsr_q(63) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(25) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(55) xor data_in(56) xor data_in(58) xor data_in(59) xor data_in(61) xor data_in(63);
    lfsr_c(29) <= lfsr_q(0) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(25) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(36) xor lfsr_q(41) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(53) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(62) xor lfsr_q(63) xor data_in(0) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(25) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(36) xor data_in(41) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(50) xor data_in(51) xor data_in(53) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(62) xor data_in(63);
    lfsr_c(30) <= lfsr_q(1) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(26) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(42) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(54) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(63) xor data_in(1) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(26) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(37) xor data_in(42) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(49) xor data_in(51) xor data_in(52) xor data_in(54) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(63);
    lfsr_c(31) <= lfsr_q(0) xor lfsr_q(4) xor lfsr_q(6) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(25) xor lfsr_q(26) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(51) xor lfsr_q(55) xor lfsr_q(63) xor data_in(0) xor data_in(4) xor data_in(6) xor data_in(18) xor data_in(20) xor data_in(22) xor data_in(25) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(32) xor data_in(33) xor data_in(36) xor data_in(37) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(55) xor data_in(63);
    lfsr_c(32) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(27) xor lfsr_q(29) xor lfsr_q(33) xor lfsr_q(35) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(46) xor lfsr_q(48) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(53) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(8) xor data_in(9) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(29) xor data_in(33) xor data_in(35) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(48) xor data_in(50) xor data_in(51) xor data_in(53) xor data_in(56) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(63);
    lfsr_c(33) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(30) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(41) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(50) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(61) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(8) xor data_in(10) xor data_in(13) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(21) xor data_in(30) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(41) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(50) xor data_in(53) xor data_in(54) xor data_in(57) xor data_in(58) xor data_in(61) xor data_in(63);
    lfsr_c(34) <= lfsr_q(1) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(9) xor lfsr_q(11) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(31) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(42) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(51) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(62) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(9) xor data_in(11) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(22) xor data_in(31) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(42) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(54) xor data_in(55) xor data_in(58) xor data_in(59) xor data_in(62);
    lfsr_c(35) <= lfsr_q(0) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(26) xor lfsr_q(28) xor lfsr_q(32) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(53) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(58) xor data_in(0) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(47) xor data_in(48) xor data_in(50) xor data_in(51) xor data_in(53) xor data_in(55) xor data_in(56) xor data_in(58);
    lfsr_c(36) <= lfsr_q(1) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(26) xor lfsr_q(27) xor lfsr_q(29) xor lfsr_q(33) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(54) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(59) xor data_in(1) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(27) xor data_in(29) xor data_in(33) xor data_in(35) xor data_in(36) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(48) xor data_in(49) xor data_in(51) xor data_in(52) xor data_in(54) xor data_in(56) xor data_in(57) xor data_in(59);
    lfsr_c(37) <= lfsr_q(0) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(24) xor lfsr_q(27) xor lfsr_q(30) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(38) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(51) xor lfsr_q(55) xor lfsr_q(57) xor lfsr_q(59) xor lfsr_q(63) xor data_in(0) xor data_in(4) xor data_in(5) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(24) xor data_in(27) xor data_in(30) xor data_in(35) xor data_in(36) xor data_in(38) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(51) xor data_in(55) xor data_in(57) xor data_in(59) xor data_in(63);
    lfsr_c(38) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(18) xor lfsr_q(22) xor lfsr_q(24) xor lfsr_q(26) xor lfsr_q(31) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(47) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(53) xor lfsr_q(56) xor lfsr_q(59) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(18) xor data_in(22) xor data_in(24) xor data_in(26) xor data_in(31) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(38) xor data_in(39) xor data_in(41) xor data_in(42) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(53) xor data_in(56) xor data_in(59) xor data_in(63);
    lfsr_c(39) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(26) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(32) xor lfsr_q(34) xor lfsr_q(36) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(45) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(16) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(32) xor data_in(34) xor data_in(36) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(43) xor data_in(45) xor data_in(48) xor data_in(49) xor data_in(53) xor data_in(54) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(63);
    lfsr_c(40) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(12) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(26) xor lfsr_q(27) xor lfsr_q(29) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(44) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(5) xor data_in(7) xor data_in(9) xor data_in(12) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(26) xor data_in(27) xor data_in(29) xor data_in(33) xor data_in(34) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(44) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(63);
    lfsr_c(41) <= lfsr_q(1) xor lfsr_q(2) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(30) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(45) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(56) xor data_in(1) xor data_in(2) xor data_in(6) xor data_in(8) xor data_in(10) xor data_in(13) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(27) xor data_in(28) xor data_in(30) xor data_in(34) xor data_in(35) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(45) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56);
    lfsr_c(42) <= lfsr_q(2) xor lfsr_q(3) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(11) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(31) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(46) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(57) xor data_in(2) xor data_in(3) xor data_in(7) xor data_in(9) xor data_in(11) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(35) xor data_in(36) xor data_in(40) xor data_in(41) xor data_in(42) xor data_in(46) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57);
    lfsr_c(43) <= lfsr_q(3) xor lfsr_q(4) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(12) xor lfsr_q(15) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(32) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(47) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor data_in(3) xor data_in(4) xor data_in(8) xor data_in(10) xor data_in(12) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(24) xor data_in(25) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(36) xor data_in(37) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(47) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58);
    lfsr_c(44) <= lfsr_q(4) xor lfsr_q(5) xor lfsr_q(9) xor lfsr_q(11) xor lfsr_q(13) xor lfsr_q(16) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(25) xor lfsr_q(26) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(33) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(48) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor data_in(4) xor data_in(5) xor data_in(9) xor data_in(11) xor data_in(13) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(25) xor data_in(26) xor data_in(30) xor data_in(31) xor data_in(33) xor data_in(37) xor data_in(38) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(48) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(59);
    lfsr_c(45) <= lfsr_q(0) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(25) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(63) xor data_in(0) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(16) xor data_in(17) xor data_in(20) xor data_in(22) xor data_in(25) xor data_in(27) xor data_in(28) xor data_in(31) xor data_in(32) xor data_in(35) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(56) xor data_in(57) xor data_in(63);
    lfsr_c(46) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(29) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(47) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(54) xor lfsr_q(57) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(10) xor data_in(11) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(29) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(40) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(47) xor data_in(49) xor data_in(50) xor data_in(54) xor data_in(57) xor data_in(59) xor data_in(60) xor data_in(63);
    lfsr_c(47) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(3) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(28) xor lfsr_q(30) xor lfsr_q(33) xor lfsr_q(36) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(55) xor lfsr_q(59) xor lfsr_q(61) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(5) xor data_in(7) xor data_in(9) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(28) xor data_in(30) xor data_in(33) xor data_in(36) xor data_in(44) xor data_in(45) xor data_in(48) xor data_in(49) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(59) xor data_in(61) xor data_in(63);
    lfsr_c(48) <= lfsr_q(1) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(29) xor lfsr_q(31) xor lfsr_q(34) xor lfsr_q(37) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(56) xor lfsr_q(60) xor lfsr_q(62) xor data_in(1) xor data_in(2) xor data_in(4) xor data_in(6) xor data_in(8) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(29) xor data_in(31) xor data_in(34) xor data_in(37) xor data_in(45) xor data_in(46) xor data_in(49) xor data_in(50) xor data_in(53) xor data_in(54) xor data_in(56) xor data_in(60) xor data_in(62);
    lfsr_c(49) <= lfsr_q(2) xor lfsr_q(3) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(11) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(30) xor lfsr_q(32) xor lfsr_q(35) xor lfsr_q(38) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(57) xor lfsr_q(61) xor lfsr_q(63) xor data_in(2) xor data_in(3) xor data_in(5) xor data_in(7) xor data_in(9) xor data_in(11) xor data_in(13) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(30) xor data_in(32) xor data_in(35) xor data_in(38) xor data_in(46) xor data_in(47) xor data_in(50) xor data_in(51) xor data_in(54) xor data_in(55) xor data_in(57) xor data_in(61) xor data_in(63);
    lfsr_c(50) <= lfsr_q(3) xor lfsr_q(4) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(12) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(31) xor lfsr_q(33) xor lfsr_q(36) xor lfsr_q(39) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(62) xor data_in(3) xor data_in(4) xor data_in(6) xor data_in(8) xor data_in(10) xor data_in(12) xor data_in(14) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(24) xor data_in(31) xor data_in(33) xor data_in(36) xor data_in(39) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(52) xor data_in(55) xor data_in(56) xor data_in(58) xor data_in(62);
    lfsr_c(51) <= lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(11) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(32) xor lfsr_q(34) xor lfsr_q(37) xor lfsr_q(40) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(59) xor lfsr_q(63) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(9) xor data_in(11) xor data_in(13) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(24) xor data_in(25) xor data_in(32) xor data_in(34) xor data_in(37) xor data_in(40) xor data_in(48) xor data_in(49) xor data_in(52) xor data_in(53) xor data_in(56) xor data_in(57) xor data_in(59) xor data_in(63);
    lfsr_c(52) <= lfsr_q(0) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(28) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(37) xor lfsr_q(42) xor lfsr_q(46) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(54) xor lfsr_q(57) xor lfsr_q(59) xor lfsr_q(63) xor data_in(0) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(12) xor data_in(13) xor data_in(17) xor data_in(18) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(28) xor data_in(33) xor data_in(34) xor data_in(37) xor data_in(42) xor data_in(46) xor data_in(51) xor data_in(52) xor data_in(54) xor data_in(57) xor data_in(59) xor data_in(63);
    lfsr_c(53) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(2) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(16) xor lfsr_q(18) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(26) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(37) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(55) xor lfsr_q(59) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(2) xor data_in(3) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(16) xor data_in(18) xor data_in(21) xor data_in(23) xor data_in(26) xor data_in(28) xor data_in(29) xor data_in(37) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(46) xor data_in(47) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(55) xor data_in(59) xor data_in(63);
    lfsr_c(54) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(3) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(25) xor lfsr_q(26) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(53) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(3) xor data_in(5) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(14) xor data_in(16) xor data_in(17) xor data_in(21) xor data_in(22) xor data_in(25) xor data_in(26) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(34) xor data_in(35) xor data_in(37) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(49) xor data_in(53) xor data_in(56) xor data_in(58) xor data_in(59) xor data_in(63);
    lfsr_c(55) <= lfsr_q(0) xor lfsr_q(1) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(27) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(34) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(41) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(63) xor data_in(0) xor data_in(1) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(15) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(34) xor data_in(36) xor data_in(37) xor data_in(41) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(57) xor data_in(58) xor data_in(63);
    lfsr_c(56) <= lfsr_q(1) xor lfsr_q(2) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(26) xor lfsr_q(28) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(35) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(42) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(58) xor lfsr_q(59) xor data_in(1) xor data_in(2) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(13) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(26) xor data_in(28) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(35) xor data_in(37) xor data_in(38) xor data_in(42) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(48) xor data_in(49) xor data_in(52) xor data_in(53) xor data_in(54) xor data_in(55) xor data_in(58) xor data_in(59);
    lfsr_c(57) <= lfsr_q(0) xor lfsr_q(3) xor lfsr_q(4) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(16) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(23) xor lfsr_q(27) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(63) xor data_in(0) xor data_in(3) xor data_in(4) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(11) xor data_in(12) xor data_in(16) xor data_in(17) xor data_in(18) xor data_in(20) xor data_in(23) xor data_in(27) xor data_in(28) xor data_in(29) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(39) xor data_in(41) xor data_in(42) xor data_in(43) xor data_in(47) xor data_in(48) xor data_in(51) xor data_in(52) xor data_in(54) xor data_in(55) xor data_in(56) xor data_in(58) xor data_in(63);
    lfsr_c(58) <= lfsr_q(1) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(17) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(21) xor lfsr_q(24) xor lfsr_q(28) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(52) xor lfsr_q(53) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(59) xor data_in(1) xor data_in(4) xor data_in(5) xor data_in(7) xor data_in(8) xor data_in(9) xor data_in(12) xor data_in(13) xor data_in(17) xor data_in(18) xor data_in(19) xor data_in(21) xor data_in(24) xor data_in(28) xor data_in(29) xor data_in(30) xor data_in(32) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(40) xor data_in(42) xor data_in(43) xor data_in(44) xor data_in(48) xor data_in(49) xor data_in(52) xor data_in(53) xor data_in(55) xor data_in(56) xor data_in(57) xor data_in(59);
    lfsr_c(59) <= lfsr_q(2) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(8) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(13) xor lfsr_q(14) xor lfsr_q(18) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(22) xor lfsr_q(25) xor lfsr_q(29) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(53) xor lfsr_q(54) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(60) xor data_in(2) xor data_in(5) xor data_in(6) xor data_in(8) xor data_in(9) xor data_in(10) xor data_in(13) xor data_in(14) xor data_in(18) xor data_in(19) xor data_in(20) xor data_in(22) xor data_in(25) xor data_in(29) xor data_in(30) xor data_in(31) xor data_in(33) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(41) xor data_in(43) xor data_in(44) xor data_in(45) xor data_in(49) xor data_in(50) xor data_in(53) xor data_in(54) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(60);
    lfsr_c(60) <= lfsr_q(3) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(9) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(14) xor lfsr_q(15) xor lfsr_q(19) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(23) xor lfsr_q(26) xor lfsr_q(30) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(34) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(42) xor lfsr_q(44) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(54) xor lfsr_q(55) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(61) xor data_in(3) xor data_in(6) xor data_in(7) xor data_in(9) xor data_in(10) xor data_in(11) xor data_in(14) xor data_in(15) xor data_in(19) xor data_in(20) xor data_in(21) xor data_in(23) xor data_in(26) xor data_in(30) xor data_in(31) xor data_in(32) xor data_in(34) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(42) xor data_in(44) xor data_in(45) xor data_in(46) xor data_in(50) xor data_in(51) xor data_in(54) xor data_in(55) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(61);
    lfsr_c(61) <= lfsr_q(4) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(10) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(15) xor lfsr_q(16) xor lfsr_q(20) xor lfsr_q(21) xor lfsr_q(22) xor lfsr_q(24) xor lfsr_q(27) xor lfsr_q(31) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(38) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(43) xor lfsr_q(45) xor lfsr_q(46) xor lfsr_q(47) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(55) xor lfsr_q(56) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(60) xor lfsr_q(62) xor data_in(4) xor data_in(7) xor data_in(8) xor data_in(10) xor data_in(11) xor data_in(12) xor data_in(15) xor data_in(16) xor data_in(20) xor data_in(21) xor data_in(22) xor data_in(24) xor data_in(27) xor data_in(31) xor data_in(32) xor data_in(33) xor data_in(35) xor data_in(36) xor data_in(37) xor data_in(38) xor data_in(39) xor data_in(40) xor data_in(41) xor data_in(43) xor data_in(45) xor data_in(46) xor data_in(47) xor data_in(51) xor data_in(52) xor data_in(55) xor data_in(56) xor data_in(58) xor data_in(59) xor data_in(60) xor data_in(62);
    lfsr_c(62) <= lfsr_q(0) xor lfsr_q(2) xor lfsr_q(4) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(11) xor lfsr_q(12) xor lfsr_q(14) xor lfsr_q(17) xor lfsr_q(19) xor lfsr_q(22) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(26) xor lfsr_q(32) xor lfsr_q(33) xor lfsr_q(35) xor lfsr_q(36) xor lfsr_q(39) xor lfsr_q(40) xor lfsr_q(44) xor lfsr_q(47) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(56) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(61) xor data_in(0) xor data_in(2) xor data_in(4) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(11) xor data_in(12) xor data_in(14) xor data_in(17) xor data_in(19) xor data_in(22) xor data_in(23) xor data_in(24) xor data_in(26) xor data_in(32) xor data_in(33) xor data_in(35) xor data_in(36) xor data_in(39) xor data_in(40) xor data_in(44) xor data_in(47) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(56) xor data_in(57) xor data_in(58) xor data_in(61);
    lfsr_c(63) <= lfsr_q(1) xor lfsr_q(3) xor lfsr_q(5) xor lfsr_q(6) xor lfsr_q(7) xor lfsr_q(8) xor lfsr_q(12) xor lfsr_q(13) xor lfsr_q(15) xor lfsr_q(18) xor lfsr_q(20) xor lfsr_q(23) xor lfsr_q(24) xor lfsr_q(25) xor lfsr_q(27) xor lfsr_q(33) xor lfsr_q(34) xor lfsr_q(36) xor lfsr_q(37) xor lfsr_q(40) xor lfsr_q(41) xor lfsr_q(45) xor lfsr_q(48) xor lfsr_q(49) xor lfsr_q(50) xor lfsr_q(51) xor lfsr_q(52) xor lfsr_q(57) xor lfsr_q(58) xor lfsr_q(59) xor lfsr_q(62) xor data_in(1) xor data_in(3) xor data_in(5) xor data_in(6) xor data_in(7) xor data_in(8) xor data_in(12) xor data_in(13) xor data_in(15) xor data_in(18) xor data_in(20) xor data_in(23) xor data_in(24) xor data_in(25) xor data_in(27) xor data_in(33) xor data_in(34) xor data_in(36) xor data_in(37) xor data_in(40) xor data_in(41) xor data_in(45) xor data_in(48) xor data_in(49) xor data_in(50) xor data_in(51) xor data_in(52) xor data_in(57) xor data_in(58) xor data_in(59) xor data_in(62);


    process (clk) begin
      if (clk'EVENT and clk = '1') then
        if (rst = '1') then
          lfsr_q <= b"1111111111111111111111111111111111111111111111111111111111111111";
        elsif (crc_en = '1') then
          lfsr_q <= lfsr_c;
        end if;
      end if;
    end process;
end architecture Behavioral;
